netcdf mbnrg_3b_A1B3C1D2_E1F2_E1F2_fit {
  // global attributes 
  :name = " mbnrg_3b_A1B3C1D2_E1F2_E1F2_fit";
  :k_x_intra_A_B_1 =  2.670808427321614e+00; // A^(-1))
  :k_x_intra_A_C_1 =  7.359465753687238e-01; // A^(-1))
  :k_x_intra_A_D_1 =  6.844006046514541e+00; // A^(-1))
  :k_x_inter_A_E_0 =  3.644609443422696e-01; // A^(-1))
  :k_x_inter_A_F_0 =  6.463638438491650e-01; // A^(-1))
  :k_x_intra_B_B_1 =  1.825358931225242e-01; // A^(-1))
  :k_x_intra_B_C_1 =  5.205345831907218e+00; // A^(-1))
  :k_x_intra_B_D_1 =  9.913234800555532e-01; // A^(-1))
  :k_x_inter_B_E_0 =  1.247314670847626e+00; // A^(-1))
  :k_x_inter_B_F_0 =  2.011299119161878e-01; // A^(-1))
  :k_x_intra_C_D_1 =  2.373630272318783e+00; // A^(-1))
  :k_x_inter_C_E_0 =  4.207714234102016e-01; // A^(-1))
  :k_x_inter_C_F_0 =  8.516144071301313e-01; // A^(-1))
  :k_x_intra_D_D_1 =  1.748722971242893e+00; // A^(-1))
  :k_x_inter_D_E_0 =  1.015571576525206e+00; // A^(-1))
  :k_x_inter_D_F_0 =  3.500586206828221e-01; // A^(-1))
  :k_x_intra_E_F_1 =  5.456280485350433e-01; // A^(-1))
  :k_x_inter_E_E_0 =  6.795736856613090e-01; // A^(-1))
  :k_x_inter_E_F_0 =  1.217029797021086e+00; // A^(-1))
  :k_x_intra_F_F_1 =  3.385721214231180e-01; // A^(-1))
  :k_x_inter_F_F_0 =  4.523340187415250e-01; // A^(-1))
  :ri =  4.500000000000000e+00; // A
  :ro =  5.500000000000000e+00; // A
  dimensions:
  poly = 1669;
  variables:
    double poly(poly);
data:
poly =
-7.112860490767345e+00, // 0
 2.502688322168444e+01, // 1
-8.557047642284195e+00, // 2
 1.163799456605192e+01, // 3
 1.823931565922074e+00, // 4
 4.586581856131587e+01, // 5
-2.878774819843313e+01, // 6
-2.850441544195123e+01, // 7
 1.871219339235855e+01, // 8
 2.765027841527561e+01, // 9
 3.880655264756776e+00, // 10
 7.925253888244434e+01, // 11
-7.789407937729048e+01, // 12
-3.813460485401763e+00, // 13
 2.433304189004415e+01, // 14
 2.938208299064685e+01, // 15
 1.679311872882453e+01, // 16
-7.743985610751777e+00, // 17
 3.200602158364673e+01, // 18
-1.270038497905953e+01, // 19
 5.249612854195462e+01, // 20
 4.467525716713070e+01, // 21
-5.066763297343708e+01, // 22
-3.379965615781857e+01, // 23
-7.859556042996397e+01, // 24
 5.117650379761645e+01, // 25
 7.281722063347327e+01, // 26
 1.255050934003009e+02, // 27
 3.018512614945916e+01, // 28
 1.808264897060762e+01, // 29
-6.282506002722900e+00, // 30
 3.462441332900742e+01, // 31
 5.704744356729197e+00, // 32
-1.045023646829425e+00, // 33
-4.848554453909296e+01, // 34
-5.198671303245419e+00, // 35
 2.420319786933679e+01, // 36
 4.707645762606589e-01, // 37
 1.265828873422483e+01, // 38
 1.955922409977622e+01, // 39
-2.914987444383257e+01, // 40
 8.113069007414179e+00, // 41
 2.022142035572173e+01, // 42
-8.113071280116992e+01, // 43
 9.847615436389796e-01, // 44
 2.449376957695564e+00, // 45
-2.475510626144985e+00, // 46
 1.273853185204540e+00, // 47
-1.266715163166671e+01, // 48
-3.653650792054540e+01, // 49
 1.495684925003103e+01, // 50
 4.131835311179196e+01, // 51
 4.034636909514571e+00, // 52
-9.022037300442229e+00, // 53
 4.616138263331312e+01, // 54
-1.523030589977142e+00, // 55
 8.228848309959789e+00, // 56
-1.662599881602102e+00, // 57
 9.363946652937193e+00, // 58
-5.275752219204751e+00, // 59
-2.978925272802528e+00, // 60
-2.587479847644488e+01, // 61
 1.631157956523914e+01, // 62
 3.635251616830029e+00, // 63
-6.914064004346574e+00, // 64
-1.150269990696764e+01, // 65
 9.537774560520932e+00, // 66
-3.625977544736965e+01, // 67
 1.288186057871464e+01, // 68
 1.391026978619325e+01, // 69
 3.377687617514957e+01, // 70
 1.843412916028777e+01, // 71
-2.651103064899675e+01, // 72
-4.620471939574111e+01, // 73
-7.851746287234041e+00, // 74
-1.137271209418473e+01, // 75
-3.140509578185505e+01, // 76
-3.729500540171169e+01, // 77
 1.339719049897086e+01, // 78
 2.088397914708182e+00, // 79
-1.497299762177062e+02, // 80
-5.043670487001815e+00, // 81
 9.686733744028235e+00, // 82
-5.967425480381369e+00, // 83
-5.580147847092560e+01, // 84
-2.997500608823211e+01, // 85
-1.230755822268132e+02, // 86
 1.192531909441126e+02, // 87
 4.087186348094221e+00, // 88
-7.687922835196017e+01, // 89
 5.788950103622580e+00, // 90
-1.157037421374161e+01, // 91
-8.533279696457811e+01, // 92
 1.822058651604981e+02, // 93
-1.443299719455538e+02, // 94
 3.815465867194974e+01, // 95
 5.482481550542068e+01, // 96
-6.770913859281930e+01, // 97
-2.854708747707874e+01, // 98
 1.508274183685035e+00, // 99
-1.488968815450214e+02, // 100
-4.782904052391665e+01, // 101
 1.415251097037149e+01, // 102
-1.258640166692962e+02, // 103
-1.114066616167136e+02, // 104
 4.439906952455411e+01, // 105
 6.694175508310343e+01, // 106
-3.814591267713401e+01, // 107
 2.646426522427549e+01, // 108
-2.577495695791394e+01, // 109
 2.324693426818179e+01, // 110
 2.350129341456957e+01, // 111
-5.170433840393110e+01, // 112
-8.796007752699753e+00, // 113
-1.566385321894453e-01, // 114
 8.234961613420511e+00, // 115
 1.419903690479060e+02, // 116
-2.420770372955004e+02, // 117
-4.861327992645534e+01, // 118
-5.305547760033175e+00, // 119
 2.572012775438875e+01, // 120
 2.850281514424068e+01, // 121
-1.071449688806481e+02, // 122
 3.868671084123019e+01, // 123
-3.213127950480359e+01, // 124
-4.490730359855764e+01, // 125
 5.027474468381078e+01, // 126
-1.168967382898540e+02, // 127
-6.982995361319382e+01, // 128
-2.394202560724675e+02, // 129
-6.176618405578071e+00, // 130
 1.016168277022537e+00, // 131
-1.411476266258695e+02, // 132
-7.939892972306394e+01, // 133
 1.484651303535035e+02, // 134
 3.669198243040057e+01, // 135
-1.478565385157064e+02, // 136
 8.054602146478342e+01, // 137
-1.119709307385752e+02, // 138
-2.589639353383874e+01, // 139
-5.260624131675994e+01, // 140
-1.319201442299155e+01, // 141
 2.302872928429375e+01, // 142
 5.866691395898940e+01, // 143
 9.107040249660955e+00, // 144
-7.356156638354918e+01, // 145
-1.297335658247520e+01, // 146
-1.659367095192275e+01, // 147
 6.689553772354284e+01, // 148
 2.998914637126710e+01, // 149
 5.066086959438608e+01, // 150
 2.907082526044476e+01, // 151
-4.908496811366855e+01, // 152
 1.605320795839703e+01, // 153
-8.122446145656173e+00, // 154
 5.104661504114981e+01, // 155
-3.752188793235474e+01, // 156
 1.636019349795129e+01, // 157
-1.170738539941569e+02, // 158
-1.765008111805632e+02, // 159
-7.988290361083703e+01, // 160
-9.867577083817058e-01, // 161
 2.061708910643641e+00, // 162
-7.167731764580029e+01, // 163
 3.564829961797810e+01, // 164
-2.210735604387015e+01, // 165
 2.719827890714524e+01, // 166
-2.690920742520801e+01, // 167
 1.634206953825526e+01, // 168
 4.147875315190646e+01, // 169
-4.650948560670781e+01, // 170
-1.975381443390921e+01, // 171
 1.649070019918317e+01, // 172
 3.550412635592854e+00, // 173
 8.949283784777541e-01, // 174
 5.791065402315240e+01, // 175
 1.024948918541486e+02, // 176
-5.241549707834562e+00, // 177
 1.027018671885152e+00, // 178
 2.572799130590762e+01, // 179
 3.124261322541789e+01, // 180
-1.081563346619756e+02, // 181
-5.158727947366796e+01, // 182
 9.578892084029889e+00, // 183
-1.521437922546390e+02, // 184
-2.758705604962318e+02, // 185
 4.145135316651336e+01, // 186
-1.360612201852886e+00, // 187
 1.135555007002180e+02, // 188
 1.845798857172833e+01, // 189
-7.993409842236909e+01, // 190
 1.399639418582152e+01, // 191
 7.322639964797972e+01, // 192
 4.134826877196270e+00, // 193
-7.394831575005257e+01, // 194
 5.527369480007868e+01, // 195
-6.486948205664218e+01, // 196
-8.370969328044798e+01, // 197
-4.585791831900794e+01, // 198
 7.751059026592161e+01, // 199
 1.122924396816331e+02, // 200
 6.845783173534126e+00, // 201
 4.383604387699237e+01, // 202
-3.722234788991964e+01, // 203
-1.581537840641696e+01, // 204
 4.563663265954311e+01, // 205
 1.411498085503614e+01, // 206
-1.006927099217001e+02, // 207
 8.493005782770732e+01, // 208
 5.465316501806777e+01, // 209
-2.105237031673123e+01, // 210
 4.901508648968368e+00, // 211
 2.096690869353950e+01, // 212
-2.507979607540325e+01, // 213
-1.675759145394714e+01, // 214
 1.702939243454925e+01, // 215
-5.467538911601462e+01, // 216
 1.554694691410176e+01, // 217
 5.666291447207129e+01, // 218
 1.386498248773010e+02, // 219
 1.663315668924014e+01, // 220
 1.336021690536708e+01, // 221
 5.106892473678059e+00, // 222
-1.919675638944354e+01, // 223
-8.118922016638992e+01, // 224
 2.009787082472758e+01, // 225
 1.374741599350302e+02, // 226
-1.249712029591604e+01, // 227
-1.191531969702133e+01, // 228
-8.513749130291950e+00, // 229
-1.277764468603102e+02, // 230
-9.362289590158416e+01, // 231
-1.590052793235282e+02, // 232
-5.920817086159975e+01, // 233
-2.911790786043237e+01, // 234
 8.163335943109804e+00, // 235
 7.234558198458154e+01, // 236
 1.748151262200398e+01, // 237
-2.874263015664216e+01, // 238
-1.731665864645214e+01, // 239
 1.913121063330907e+01, // 240
 1.220759038571246e+01, // 241
 2.266890159535852e+00, // 242
 4.960933001188685e+00, // 243
-1.848303800938552e+01, // 244
 1.959388665249793e+02, // 245
 1.490173241606080e+01, // 246
 1.665658505197978e+01, // 247
-8.162151792391005e-01, // 248
-3.180309944787875e+01, // 249
-1.195159317499606e+01, // 250
 2.858214826134539e+01, // 251
-1.559455271210255e+02, // 252
-1.541312164861104e+01, // 253
-2.557070404318381e+01, // 254
-3.175714216535686e+00, // 255
 8.371600791278792e+01, // 256
-6.022740057013743e+01, // 257
 3.140932081273429e+01, // 258
 1.372165490917584e+02, // 259
-1.008393225091754e+01, // 260
-1.158397719815370e+02, // 261
-1.266956536322142e+01, // 262
-3.490994951220322e+01, // 263
-1.563936793854185e+01, // 264
 1.836995621552238e+02, // 265
-3.916639040376893e+01, // 266
-2.128273949088343e+01, // 267
 3.264828462160848e+00, // 268
 3.431523145849908e+01, // 269
-7.900743078808062e-01, // 270
 1.168362873311881e+02, // 271
 9.168489972586664e-01, // 272
-1.094929216839270e+02, // 273
 4.638781147201169e+01, // 274
 3.052719368988927e+01, // 275
-2.943670907481053e+01, // 276
 2.937411113136980e+01, // 277
-1.375609640055098e+01, // 278
-1.503667336313328e+02, // 279
 4.667482251971470e+01, // 280
 2.713597237366292e+01, // 281
-9.039654064652089e+01, // 282
 4.332057163341635e+01, // 283
-1.696217265947548e+02, // 284
-1.300523911105101e+02, // 285
 2.576584613382449e+00, // 286
-2.231190900144765e+01, // 287
 3.555431673185966e+01, // 288
 7.171443404798919e+01, // 289
 8.868230336593729e-01, // 290
-1.143874777469002e+02, // 291
-3.121467285509899e+01, // 292
-9.736171327980824e+01, // 293
 1.858120344317006e+01, // 294
-4.105975833168587e+01, // 295
 6.102216897741735e+01, // 296
 8.153015107724107e+01, // 297
-2.917696997686258e+01, // 298
-2.850421356152525e+00, // 299
 5.572411587921281e+00, // 300
-1.600714539979367e+02, // 301
-3.043417799829308e+01, // 302
 9.492275574875778e+01, // 303
-1.431451976355915e+02, // 304
 2.573732845052712e+00, // 305
-1.651079136984114e+01, // 306
 2.719475859223744e+01, // 307
-5.322339363305038e+01, // 308
 4.911925171606445e+01, // 309
-3.218253266388327e+01, // 310
-2.662912679881797e+01, // 311
 2.748206731828148e+00, // 312
 7.000062886447250e+01, // 313
-1.853096144171804e+01, // 314
-2.936792119967998e+01, // 315
 1.481558080558231e+01, // 316
-2.116439008837531e+01, // 317
-8.622335567437737e+00, // 318
 3.522814142648266e+01, // 319
-2.563248339755760e+01, // 320
 2.479775987967599e+01, // 321
-2.215233849331878e+01, // 322
-9.226403316950096e+01, // 323
-3.668222772654151e+01, // 324
 1.361127744837727e+01, // 325
-2.215717418715713e+01, // 326
 1.302166641574499e+02, // 327
 4.124651088807501e+00, // 328
-4.176292330328825e+01, // 329
-2.158184567610084e+01, // 330
 8.150763661464836e+01, // 331
 1.008455746995575e+02, // 332
-8.592910584620442e+01, // 333
 5.311258823601743e+01, // 334
 1.212198977936378e+02, // 335
-2.583081024689083e+00, // 336
-3.180427026075796e+01, // 337
 1.204621161320661e+01, // 338
 3.904469141112695e+00, // 339
-9.706250711965224e+01, // 340
 1.166806277045581e+01, // 341
 1.523459646752172e+02, // 342
-1.893913915976685e+01, // 343
 4.849531268813351e+00, // 344
-4.816789107769203e+00, // 345
 6.783075394935054e+01, // 346
 1.308459142609425e+01, // 347
-1.166403854485119e+02, // 348
-8.051282203833571e+00, // 349
 4.564361543586950e+00, // 350
-8.819349737294836e+00, // 351
 1.915896721757124e+01, // 352
 6.081278729237105e+01, // 353
 2.050586370597984e+00, // 354
 2.117918172969296e+00, // 355
 2.511559729461034e+01, // 356
-1.967850194518307e+01, // 357
-8.875136833419153e+01, // 358
 6.288373927087345e+01, // 359
-1.448274221695999e+01, // 360
 1.187095908836710e+01, // 361
 7.974891025034292e+01, // 362
-1.271328087879930e+02, // 363
 4.857195695542145e+00, // 364
 3.523899836519752e+01, // 365
-5.173617548289640e+01, // 366
 1.446391919509095e+02, // 367
 9.099920384028220e+00, // 368
-1.308387965053660e+02, // 369
 7.448761298929885e+01, // 370
 2.184838258091911e+01, // 371
-1.735275803515865e+02, // 372
-1.902471513774595e+02, // 373
 4.599073165614537e+00, // 374
 3.232031152462539e+01, // 375
-3.432259182441657e+01, // 376
-1.701601919604460e+01, // 377
-2.042843588927760e+02, // 378
-1.023296207896284e+01, // 379
-7.632125677084689e+01, // 380
-5.595311335529045e+01, // 381
 7.152451601293592e+01, // 382
-1.526597097909621e+02, // 383
 7.971038780446031e+01, // 384
-1.453992952763381e+01, // 385
 1.118530736004718e+02, // 386
 4.332830438469012e-01, // 387
 4.115732058685708e+00, // 388
-2.875437442051317e+00, // 389
 1.121283514839963e+01, // 390
 1.415928798284869e+01, // 391
-1.214290349746729e+01, // 392
-2.916743809885325e+01, // 393
-2.668199580621182e+00, // 394
-3.650974493445235e+00, // 395
-2.880498782036845e+01, // 396
-1.308112128379100e+01, // 397
 6.400061172588009e-01, // 398
 4.740354972414199e+00, // 399
 3.503246796439541e+01, // 400
-1.058141404157464e+01, // 401
-3.178953817488564e+00, // 402
 9.962692747946891e+00, // 403
-2.266592051136941e+00, // 404
-2.327041111623226e+00, // 405
 8.869077905917339e-01, // 406
 3.461445966221896e+00, // 407
 1.141569382747187e-01, // 408
 8.025714925938802e+00, // 409
-3.487681266242202e+00, // 410
 1.179868903298867e+00, // 411
 2.314328874028588e+01, // 412
-1.099036594063409e+00, // 413
 1.322320875240678e+01, // 414
 2.077105431950145e+01, // 415
-1.805236818647359e+01, // 416
-1.100903359482699e+01, // 417
 3.708033564589952e+01, // 418
-2.556963240055913e+00, // 419
 2.537507016143977e+00, // 420
-2.645835740605166e+01, // 421
-3.537772632665363e+00, // 422
 1.845894567925906e+00, // 423
 2.362995571618625e+01, // 424
-2.750099352652130e+00, // 425
 6.952400628755241e+00, // 426
 8.066035573799669e+00, // 427
-1.077394238277536e+00, // 428
-9.125658881424348e-01, // 429
-1.492056403329525e+01, // 430
 5.937560482045555e+00, // 431
 3.587894683335448e+01, // 432
-3.050277245966593e+01, // 433
-1.674534737951667e+01, // 434
 8.514195820989022e+00, // 435
-9.065703131355669e+00, // 436
 5.220767533712305e+00, // 437
 2.654988357383448e+01, // 438
-1.035159217838354e+01, // 439
-3.161907796571023e+01, // 440
 2.040910913913055e+01, // 441
 3.882245284793506e-02, // 442
 9.042287532154717e+00, // 443
-4.424701921109593e+01, // 444
-8.704295703561525e+01, // 445
-8.560585533193644e+01, // 446
 6.842736249352662e+01, // 447
 4.806995082791781e+01, // 448
 7.425776822215943e+01, // 449
-1.544336222773483e+01, // 450
 4.592580439763768e+00, // 451
-9.399867548961979e+00, // 452
 1.522057452600722e+00, // 453
 4.195656886824710e+00, // 454
-9.003235209699106e-01, // 455
-7.789373274980622e+01, // 456
 1.821940423083479e+01, // 457
-9.466848173319461e-01, // 458
 1.203957128975616e+01, // 459
 1.711879595823043e+01, // 460
 8.796748946438504e+00, // 461
 2.576699309579411e+00, // 462
-5.114940919316997e+00, // 463
 4.195117603920277e+00, // 464
-3.829007048558883e+00, // 465
 3.996078242205254e+00, // 466
-2.097329233915270e+01, // 467
-7.074118891186568e+00, // 468
 1.177683516587885e+01, // 469
 2.135505363143517e+01, // 470
 3.707459130476418e+01, // 471
-1.004566422644440e+01, // 472
 2.952148451524989e-01, // 473
-1.288417196407030e+01, // 474
-1.685357384450841e+01, // 475
-2.008719770626032e+01, // 476
 1.583940971699791e+00, // 477
 1.931697547837734e+00, // 478
-2.982722522896588e-01, // 479
-4.672950652376028e+01, // 480
-4.721510206682621e+01, // 481
-2.053985538067477e+01, // 482
-6.445941188096243e+01, // 483
 3.783046719776097e+01, // 484
 3.762229073855005e+01, // 485
 2.728202669979895e+01, // 486
 7.040644127573084e+01, // 487
 1.309874557466268e+01, // 488
 1.242129633219930e+01, // 489
 4.343880959535633e+00, // 490
 4.425003503690303e+01, // 491
 6.149461791477959e+01, // 492
-2.680789435741891e+00, // 493
 1.548235322644492e+02, // 494
-2.313460528901511e+01, // 495
-4.041974062520553e+01, // 496
-1.418771562226837e+01, // 497
-7.543493462069841e+01, // 498
-1.259746638431257e+02, // 499
 3.508430344060497e+01, // 500
 2.571008534049826e+01, // 501
-3.823207524752659e+01, // 502
-6.982191044821517e-01, // 503
-8.261731678613878e-01, // 504
 1.202063652367250e+02, // 505
-1.325974884844808e+02, // 506
 7.881870991948486e+01, // 507
 1.716707524870283e+02, // 508
 4.087578943235366e+00, // 509
-8.261420939191616e+01, // 510
-4.278461922216210e+01, // 511
-1.266126636092650e+02, // 512
 1.234848361714783e+02, // 513
-5.584560254562003e+01, // 514
-1.068848166750112e+02, // 515
-1.078244220207264e+01, // 516
-1.852210887310399e+00, // 517
 6.097495476199816e+01, // 518
-4.636964761824796e+01, // 519
-2.880754373731378e+01, // 520
 5.235919572351752e+00, // 521
-1.320251402919280e+01, // 522
-2.742845139335245e+01, // 523
-2.124546134270619e+01, // 524
 8.108351158786208e+01, // 525
-6.491499410713425e+00, // 526
-3.007022857586264e+01, // 527
-1.069776311579606e+02, // 528
 1.459567999495140e+02, // 529
 4.999070860747869e+01, // 530
 1.698481342880555e+01, // 531
-1.201013453947318e+01, // 532
-1.384347504349140e+02, // 533
-2.097930665351134e+01, // 534
 3.126167439672579e+01, // 535
-9.457017925745185e+01, // 536
-5.067514514971705e+01, // 537
 2.158112328311027e+01, // 538
-1.615441183815910e+01, // 539
 5.476050614257525e+01, // 540
-1.291786087740860e+01, // 541
 4.458081638364320e+01, // 542
-1.681047509795248e+01, // 543
-2.017715229434765e+01, // 544
 1.191200804348095e+01, // 545
 1.666209040392521e+01, // 546
 8.545536441638473e+01, // 547
-8.545864810091781e+01, // 548
-3.402558150658464e+01, // 549
-1.086089510548911e+01, // 550
 9.637804832556428e+01, // 551
-3.836005095547222e+01, // 552
 6.287554116833090e+01, // 553
-2.715444927331789e+01, // 554
 7.296904373150483e+00, // 555
-3.520764576657374e+01, // 556
 7.016424694705090e+01, // 557
-4.674080612167423e+00, // 558
-1.141735802252962e+02, // 559
 8.019082471633341e+01, // 560
 9.588308967444326e+01, // 561
 7.035405158431909e+01, // 562
 6.252573066659833e+00, // 563
 3.092884835773654e+01, // 564
-4.591467782924161e+01, // 565
 1.623938852258403e+02, // 566
-2.260992939293274e+01, // 567
 8.616670830595550e+01, // 568
 1.377544417707174e+01, // 569
 4.502289531357714e+01, // 570
-4.372516219552040e+01, // 571
-2.952758508386036e+00, // 572
 8.848543390020199e+00, // 573
 8.057754489407957e+01, // 574
 6.111802518799269e+01, // 575
-2.287998933341738e+00, // 576
-1.764429419394103e+01, // 577
 9.486105099276960e+00, // 578
-2.907414593785182e+01, // 579
-1.714628969776917e+01, // 580
-1.229606108938854e+01, // 581
 6.431853253909044e+01, // 582
 3.619541935195616e+00, // 583
 9.711136948363624e+00, // 584
-3.192896596439478e-01, // 585
 2.182365369550193e+01, // 586
-5.741843068913040e+01, // 587
-4.039999612546811e+01, // 588
-9.968954749795790e+01, // 589
-9.366580291476151e+00, // 590
 4.546248612608510e+01, // 591
-1.056974268284820e+01, // 592
 2.666820493686479e+01, // 593
 1.309900709768097e+01, // 594
 5.845077524790294e+01, // 595
-7.067166850595682e+01, // 596
 2.308347233096329e+01, // 597
-4.918965489205536e+01, // 598
-2.689422232662206e+00, // 599
-3.244663232921112e+00, // 600
 2.889394678491173e+01, // 601
-1.605961454336643e+00, // 602
 3.893269265719569e+01, // 603
-2.087754579162062e+01, // 604
-3.601381400869821e-01, // 605
-8.574060759234888e+00, // 606
 4.088752582324282e+00, // 607
 6.568405532055929e+00, // 608
 3.917434985933907e+00, // 609
-3.761308785613337e+00, // 610
-1.907351712871630e+00, // 611
-1.776080893937904e+01, // 612
 1.800172813074919e+01, // 613
 2.354558843045460e+01, // 614
-3.122597467648932e+00, // 615
-9.436584054044461e+00, // 616
 3.379191211258001e+01, // 617
 8.754003869478309e+01, // 618
-2.290217626205194e+00, // 619
 1.961432399364712e+00, // 620
 6.913563687253119e+00, // 621
-1.852643887685444e+01, // 622
 5.344724598735291e+01, // 623
-1.211470871574064e+01, // 624
 2.271509180859433e+01, // 625
 4.477570759213878e+00, // 626
 1.765889083491243e+01, // 627
 2.914478888069620e+00, // 628
 4.778812977692235e+01, // 629
-2.332943040185430e+01, // 630
 6.362106801945341e+00, // 631
-1.865682377423555e+00, // 632
-1.542385418352854e+00, // 633
 1.487612423165132e-01, // 634
-5.978254584900240e-01, // 635
 2.211013927260880e+01, // 636
-3.764206837502491e+01, // 637
 4.030036597772141e+01, // 638
-3.680799330135465e+01, // 639
 3.951587425837100e+00, // 640
-1.339406226288990e+01, // 641
-2.177073978726885e+00, // 642
 2.897196866588266e-01, // 643
 1.746238541182187e+01, // 644
-1.007686927833366e+02, // 645
-5.854124611998153e+01, // 646
-4.613920825089949e+01, // 647
-2.993743004320959e+01, // 648
 7.401080401451215e+00, // 649
 1.744751679647161e+01, // 650
 1.780136312465753e+01, // 651
 5.963465140105934e+00, // 652
 6.015544739078938e+00, // 653
 1.715870039953169e+01, // 654
 4.867266913425500e+01, // 655
-4.140760389441061e+01, // 656
-2.187153882051470e+00, // 657
-9.028394621224923e+00, // 658
 5.973586167688451e+00, // 659
-1.988610781181228e+01, // 660
-1.256114869236644e+01, // 661
 3.641945076573066e+00, // 662
 4.839507812449253e+00, // 663
 8.554449764150792e+00, // 664
-7.357342000890606e+01, // 665
-2.071178286616318e+01, // 666
-2.662009377052034e+01, // 667
-1.231899383359552e+01, // 668
-2.012070569651005e+01, // 669
-1.035923886712782e+01, // 670
-2.019983874817195e+00, // 671
-1.414522416587250e+01, // 672
-1.888983979616004e+01, // 673
 5.637337775018469e+01, // 674
-5.854706005728178e+01, // 675
-3.488043487521772e+01, // 676
 1.248683947689557e+01, // 677
 2.438938016966790e+00, // 678
 6.036358195317157e+00, // 679
 4.346495326979308e+00, // 680
 6.567944433743924e+01, // 681
 4.501262856909067e+01, // 682
-6.702378580891263e+00, // 683
 1.337926971838545e+01, // 684
 1.209357431070015e+01, // 685
 2.811464565977309e+00, // 686
 3.614420415570464e+00, // 687
 5.055939416410105e+00, // 688
 1.388622927892074e+00, // 689
 6.770732061704837e+00, // 690
-2.289643308617145e+01, // 691
-1.775798510304804e+01, // 692
-2.149539546645042e+01, // 693
-2.063999141481943e+01, // 694
 1.696172724573491e+00, // 695
-8.079750251624299e+00, // 696
 2.043467973179762e+01, // 697
 2.573269826159658e+01, // 698
-7.312515365655845e+00, // 699
 6.354754827545266e+01, // 700
 7.187839755862930e+00, // 701
 1.371931273065660e+01, // 702
 1.866864701417074e+01, // 703
 4.492273967941367e+01, // 704
-3.972300748198919e+01, // 705
-1.160988272625806e+01, // 706
 5.267983440703840e+01, // 707
 2.223020907478636e+01, // 708
 1.849078296186121e+01, // 709
 1.010540074630635e+02, // 710
-1.821527550258856e+01, // 711
-1.388663588823846e+01, // 712
-1.945706419581087e+01, // 713
 8.725325303960080e+00, // 714
 2.150851522740998e+01, // 715
 1.146370812898199e+01, // 716
-1.265332502405496e+01, // 717
 3.823476654783872e+01, // 718
 1.307083686236991e+01, // 719
 4.893129536234685e+01, // 720
 6.181231401359702e+01, // 721
-3.627525933529453e+00, // 722
 7.674999032813590e+00, // 723
-1.940148082768478e+01, // 724
-8.989143801622642e+00, // 725
 5.339438848538887e+01, // 726
-8.668688014018694e-01, // 727
 5.183761835355446e+01, // 728
 1.481471450731142e+01, // 729
-6.898373358699368e+01, // 730
 2.066141126056058e+01, // 731
 5.652336213937092e+01, // 732
-2.143712278409439e+01, // 733
-4.270997803092055e+01, // 734
 3.785465426746009e+01, // 735
 7.651545669069169e+00, // 736
 2.991221683404722e+01, // 737
 1.050206829594731e+02, // 738
 1.456782916583607e+02, // 739
 7.537541583827128e+01, // 740
-1.101949111559648e+02, // 741
-2.752557273387050e+01, // 742
-9.928168556042370e+01, // 743
 5.443774165869793e+01, // 744
-3.482812806949868e+01, // 745
 2.066209534973686e+01, // 746
-7.533598411517315e+01, // 747
 3.240209240767192e+01, // 748
-6.196495018424965e+01, // 749
 3.618416199873398e+01, // 750
-2.146037898529758e+01, // 751
 3.796351065320379e+01, // 752
 1.637236072632071e+01, // 753
-1.045273105166984e+01, // 754
-4.845110683329486e+01, // 755
 9.373595333983353e+01, // 756
-4.433208472405958e+01, // 757
-5.729643978099296e+01, // 758
 4.917090588887199e+01, // 759
 5.276880944856877e+01, // 760
 4.218405038505208e+00, // 761
-2.006140748048680e+01, // 762
 3.017255555972513e+01, // 763
-1.781394625440063e+01, // 764
 3.646513314229636e+01, // 765
 5.418610136790904e+01, // 766
 1.028606326538512e+01, // 767
 5.813948905951477e+00, // 768
-3.748472375377960e+01, // 769
-4.096061857550576e+00, // 770
-1.216283303544731e+02, // 771
-5.529467037989868e+01, // 772
 1.381822156644425e+02, // 773
-4.417352291586206e+01, // 774
 4.118265743877226e+01, // 775
 1.950479860535693e+01, // 776
 2.393630477073206e+01, // 777
 6.258650377460321e+01, // 778
 1.873164200853205e+01, // 779
 7.398041791941419e+01, // 780
-4.839369953839815e+01, // 781
 1.265768602696475e+01, // 782
 1.059355371763264e+02, // 783
-6.434666220753323e+01, // 784
 1.202504113599233e+01, // 785
-4.378509380988734e+01, // 786
 3.006805073242377e+01, // 787
 1.700576976632094e+02, // 788
 1.688090915340133e+01, // 789
-5.577955839670688e+01, // 790
 5.643943814552044e+01, // 791
-3.614836420792090e+01, // 792
-6.291776887507282e+00, // 793
 1.492822450459758e+01, // 794
-6.367839666721269e+00, // 795
-1.816004116515213e+01, // 796
 3.770508754379774e+01, // 797
-1.530429996489937e+01, // 798
 1.555838498692284e+01, // 799
-2.502952389046444e+01, // 800
 7.552303939724368e+01, // 801
-1.199686426584751e+01, // 802
 2.530584007147930e-01, // 803
-5.977795725775206e+01, // 804
 6.407004510727860e+00, // 805
-3.698062913518880e+01, // 806
 2.949270383953966e+01, // 807
-1.501285482528581e+01, // 808
 9.730746345253738e+00, // 809
 1.480858349864959e+01, // 810
-6.950892984651247e+00, // 811
-7.042600741827059e+01, // 812
-1.525087350448895e+01, // 813
-1.194054363429768e+02, // 814
-6.584302728072662e+01, // 815
-2.633945366797604e+01, // 816
 5.743699527704557e+01, // 817
 8.068362736306268e+01, // 818
 2.077343213674062e+01, // 819
-1.023924283974111e+01, // 820
-1.246708375554534e+01, // 821
-6.569164790714122e+00, // 822
-5.613357299744033e+00, // 823
-3.780469393273986e+01, // 824
-1.119485035497994e+02, // 825
 6.871266850457718e+01, // 826
 6.198825552463161e+01, // 827
 1.640708691207736e+01, // 828
 4.205188285926187e+01, // 829
 2.808588869702583e+01, // 830
 1.001207486220602e+00, // 831
-1.974114916298648e+01, // 832
 2.497631234178738e+01, // 833
-9.534185556685680e+00, // 834
 1.646865667916752e-02, // 835
 2.955547824144316e+01, // 836
 6.689358822764886e+01, // 837
-4.855351840822098e+01, // 838
 7.277342047285747e+00, // 839
-5.605217827507223e+00, // 840
 2.774247267982219e+01, // 841
 1.863993651176405e+01, // 842
 2.425363797626434e+01, // 843
 4.409074454776628e+01, // 844
 1.319408617723901e+01, // 845
 1.836092512115712e+00, // 846
 1.571230711613028e+01, // 847
 6.864511940249761e+00, // 848
-7.751141423135191e+01, // 849
-4.791814413401143e+01, // 850
 2.455392890589403e+01, // 851
 2.478493035002155e+00, // 852
 3.999320581094578e+01, // 853
 3.554428920486924e+01, // 854
 2.506698728495101e+01, // 855
-8.238033519018499e+01, // 856
 3.334574355957130e+01, // 857
-7.366158766151320e+01, // 858
 6.848619363618372e+00, // 859
-9.279333473143095e+01, // 860
 3.287467989980247e+01, // 861
 2.679613904057994e+01, // 862
 2.411867020232560e+00, // 863
-1.003470795927265e+00, // 864
 1.659092298659480e+01, // 865
 3.868815226600044e+01, // 866
-1.114133224882597e+01, // 867
-3.634057145529385e+01, // 868
 3.691599282560482e+01, // 869
 3.013353461810599e+01, // 870
-2.363086237506721e+00, // 871
-2.028951351040349e+01, // 872
-1.182792292405738e+01, // 873
-1.072367793926255e+02, // 874
-1.067989699555240e+02, // 875
 1.353637411645628e+00, // 876
-1.690286380874696e+01, // 877
-6.276601226094420e+01, // 878
 3.764579916948171e+01, // 879
 6.276239907342030e+01, // 880
 2.188934103464987e+01, // 881
-1.327483502646847e+01, // 882
 1.552894337907061e+02, // 883
 2.778068691142573e+01, // 884
 5.938622219884618e+00, // 885
-2.782684875242760e+01, // 886
-4.612343609778670e+01, // 887
-2.922339676786296e+01, // 888
 3.489734671204478e+01, // 889
 2.169109340373986e+01, // 890
-2.279523027084465e+01, // 891
 7.744422986937916e+00, // 892
 1.955290768016031e+02, // 893
 2.530554494834310e+01, // 894
 1.616277773982552e+01, // 895
 1.844260129630653e+01, // 896
 2.369826401945558e+01, // 897
-1.020427363415253e+02, // 898
-6.063906274783879e+01, // 899
-3.930743664740383e+01, // 900
-8.014189315031963e+00, // 901
-4.067669125017069e+00, // 902
 1.539273746663712e+01, // 903
 1.278591029636010e+02, // 904
 5.878135816355989e-01, // 905
-4.969993407091766e+01, // 906
-1.555135847747328e+01, // 907
-6.843279100271725e+01, // 908
 2.286876307719610e+01, // 909
-7.910617573469772e+00, // 910
-9.556042947294359e-02, // 911
 2.768168784129677e+01, // 912
 1.462703034691453e+01, // 913
-1.607515115946906e+01, // 914
 6.918582945886888e+01, // 915
-7.130467357642337e+00, // 916
-2.000043128089772e+01, // 917
-8.370314411484937e+01, // 918
-1.773591439296104e+01, // 919
-2.145634422868309e+01, // 920
-2.176714882223341e+01, // 921
 3.760149606683974e+01, // 922
 1.141717657799156e+02, // 923
-5.679487248816353e+01, // 924
-1.288592394405468e+02, // 925
 9.734151616851072e+01, // 926
-3.180253526756571e+01, // 927
 1.816982767445222e+01, // 928
 6.485382737579158e+01, // 929
 6.021028038800839e+01, // 930
 9.505797822597332e+01, // 931
-1.204491205694088e+02, // 932
 6.988594573847874e+01, // 933
-1.556222732921141e+01, // 934
 3.252371569584124e+01, // 935
 1.745985914534768e+01, // 936
-7.378092337975289e+01, // 937
 4.079491229183911e+01, // 938
-6.504627684890077e+00, // 939
-1.422587017321680e+01, // 940
 8.662201750590604e+00, // 941
 1.475449180921826e+00, // 942
-8.205725069825794e+00, // 943
-8.802185521529724e+01, // 944
-7.905707078848323e+00, // 945
-1.144720423694331e+01, // 946
-8.178389304188403e+00, // 947
 2.995155080314058e+01, // 948
-2.536924857014259e+01, // 949
-9.920189178360788e+00, // 950
 3.030777368704473e+01, // 951
 2.798802100554866e+01, // 952
-5.953018441228544e+00, // 953
-3.761950889201289e-01, // 954
-3.505964553163654e+01, // 955
 3.720942076258415e+01, // 956
-1.504665079915040e+01, // 957
 7.730335806369123e+01, // 958
 2.686878421605012e+01, // 959
 7.584154400631343e+01, // 960
-3.812397225197493e+00, // 961
 1.679794953962178e+01, // 962
 5.591940562493316e+00, // 963
 5.982400680259646e+01, // 964
-3.006947390490642e+01, // 965
-4.114743303291387e+01, // 966
 7.711887808270996e+00, // 967
 9.646015310177567e+01, // 968
-1.293904983591093e+01, // 969
 1.286410001348036e+02, // 970
 8.866788789230290e+00, // 971
 4.495817777895322e+01, // 972
-1.599584130795116e+01, // 973
 2.085356556670807e+01, // 974
-5.119002683605757e+00, // 975
-1.711775592621961e+01, // 976
 1.618518673955857e+01, // 977
-2.020246909374078e+01, // 978
 6.756271037440804e+01, // 979
-3.071817348270718e+01, // 980
 1.673076853072211e+02, // 981
-9.505955093521244e+00, // 982
-3.782142078136165e+01, // 983
 2.177131787582132e+00, // 984
-1.169815495634925e+02, // 985
 4.592801735997267e+00, // 986
-1.138489691861759e+02, // 987
-3.332694763208988e+01, // 988
-3.807250867578110e+01, // 989
 1.531639979030823e+00, // 990
 5.615948316178661e+01, // 991
-3.879278198063157e+01, // 992
 3.691881016083192e+01, // 993
 9.059970430415601e+01, // 994
 8.032912332220801e+01, // 995
-1.069055319616434e+02, // 996
 1.131407257195658e+02, // 997
-3.601449848473298e+01, // 998
 1.606890025211769e+01, // 999
-1.678147918846573e+01, // 1000
 3.674381310827090e+01, // 1001
 3.650202088492847e+01, // 1002
-4.852381697141021e+01, // 1003
-8.485107406850344e+01, // 1004
-5.825371274237994e+01, // 1005
-1.711182420680046e+01, // 1006
-7.264335181710595e+00, // 1007
-1.381179601258894e+02, // 1008
 2.815921996180986e+01, // 1009
 7.621652494929710e+01, // 1010
 1.144948708603344e+02, // 1011
-4.740727395201165e+00, // 1012
 4.230758028850738e+01, // 1013
 8.217072226594770e+00, // 1014
-4.611837217330986e-01, // 1015
-1.727734429058889e+01, // 1016
-7.338596437955842e+01, // 1017
 2.066098516130175e+01, // 1018
-1.398856135292472e+01, // 1019
 2.332985263169448e+01, // 1020
 7.312800520900737e+01, // 1021
 1.779083328275250e+00, // 1022
-3.260563867712228e+01, // 1023
 2.497700910756866e+02, // 1024
 6.218387838471183e+01, // 1025
 1.568399965606555e+02, // 1026
 1.196003189072200e+01, // 1027
-5.507226113511295e+01, // 1028
-7.702594232770664e+01, // 1029
 4.720610157245982e+01, // 1030
 1.151301532568963e+02, // 1031
 1.835998115688633e+01, // 1032
-2.887962018979230e+00, // 1033
-7.987032143123328e+01, // 1034
 8.945625694057655e+01, // 1035
 7.723524945192732e+01, // 1036
-2.528747543639895e+01, // 1037
 6.089290305998826e+00, // 1038
 5.964610622346330e+00, // 1039
-7.570404568622634e+01, // 1040
-8.165938523428989e+01, // 1041
-2.696603166896628e+01, // 1042
-2.512648402605085e+01, // 1043
 4.179975009769343e+01, // 1044
 1.382115065804570e+01, // 1045
-3.766783444121112e+00, // 1046
-2.998236840633074e+01, // 1047
-1.918603327339574e+01, // 1048
 3.422893686547355e+00, // 1049
-4.721252417286259e+01, // 1050
-1.409491530094549e+01, // 1051
-9.652148480776848e+00, // 1052
-1.232979760941433e+01, // 1053
 7.580081764829025e-02, // 1054
-6.897438595494157e+01, // 1055
-2.766540216556827e+01, // 1056
-9.729192945703515e+00, // 1057
-3.325899830971959e+01, // 1058
 1.359303038206976e+01, // 1059
-5.679599211622829e+01, // 1060
-1.969941052156435e+01, // 1061
 2.361350757507986e+02, // 1062
 1.248495454802841e+02, // 1063
-3.488531246708838e+01, // 1064
-1.907979571741195e+01, // 1065
 1.542258724814878e+02, // 1066
 5.715971830535187e+01, // 1067
-1.418106982333756e+02, // 1068
 2.769761017383158e+01, // 1069
-1.538938378537206e+01, // 1070
-1.509973300396711e+00, // 1071
 1.365141470414504e+02, // 1072
 9.608866036100676e+01, // 1073
-3.343737072552212e+01, // 1074
 9.575107522883663e+01, // 1075
-7.807807508771977e+01, // 1076
-9.017468988618267e+00, // 1077
 1.910694251421950e+00, // 1078
 1.000577946763545e+01, // 1079
-3.542432109022173e+01, // 1080
-9.136284813866656e+00, // 1081
-7.843343240617252e+00, // 1082
-4.183122948005946e+01, // 1083
 6.203079915998019e+00, // 1084
 1.139499785625621e+01, // 1085
 7.366486704112107e+01, // 1086
 6.616853405901546e+00, // 1087
-1.043646446745959e+00, // 1088
-2.114105754842408e+01, // 1089
 1.469045726030722e+01, // 1090
 1.981267564033059e+01, // 1091
 6.215310910604104e+00, // 1092
-5.110664575007207e+00, // 1093
-1.265009577030646e+01, // 1094
 4.845454544774029e+01, // 1095
-1.751101378874128e+01, // 1096
-2.756236448923646e+00, // 1097
-1.050650184686632e+01, // 1098
-2.616581226699155e+00, // 1099
 5.847260200744991e+00, // 1100
-9.765113346887100e-01, // 1101
 4.985570116446846e+00, // 1102
 3.504930275052958e+01, // 1103
-1.159828136180524e+01, // 1104
 2.965820635722441e+01, // 1105
 8.880312004223912e+01, // 1106
 2.422193458444491e+01, // 1107
-1.786492793716153e+01, // 1108
-7.322986279639738e+01, // 1109
-1.223371939124598e+02, // 1110
-8.524226395513037e+01, // 1111
-1.211428642630726e+02, // 1112
 2.854750407789995e+01, // 1113
-4.991569327778670e+00, // 1114
 1.710484770331185e+01, // 1115
 3.670087671163435e+01, // 1116
-6.827692474130785e+01, // 1117
-1.090465202687043e+00, // 1118
 7.692890498002619e+00, // 1119
 8.000326555131070e+01, // 1120
-8.222368924484250e+01, // 1121
 5.626363175942678e+01, // 1122
-1.393337953281915e+02, // 1123
-2.414144037921698e+00, // 1124
 1.272387196466599e+01, // 1125
 1.384489175502033e+01, // 1126
-6.918703512577650e+01, // 1127
 8.588557911538443e+00, // 1128
-2.170533260828698e+01, // 1129
 1.143015099573959e+00, // 1130
 4.677806898868671e-01, // 1131
-3.824208253832765e+01, // 1132
 1.547626447337934e+01, // 1133
 5.786935805557987e+01, // 1134
-2.236814991664759e+01, // 1135
-3.939059199927839e+01, // 1136
 4.411823430964685e+00, // 1137
 2.442785364328681e+01, // 1138
 2.375395358350619e+01, // 1139
-5.406472834771927e+00, // 1140
 1.177188006892508e+01, // 1141
-4.518492757957125e+00, // 1142
 7.510376599264999e+00, // 1143
-9.078055984630492e+00, // 1144
 1.206837497181398e+01, // 1145
-1.123824125047783e+00, // 1146
 1.180327560871743e+01, // 1147
 2.340379032540874e+01, // 1148
-3.527109102865568e+01, // 1149
-1.166019929349232e+00, // 1150
 3.723166614354385e+01, // 1151
 2.824185231701561e+00, // 1152
 1.987748493952457e+01, // 1153
 8.318827389881567e+01, // 1154
-8.563407755264852e+01, // 1155
-7.231396178346850e+00, // 1156
 3.375604266759426e+01, // 1157
-1.782946461536191e+02, // 1158
 9.051198767231803e+01, // 1159
 8.411052450468118e+01, // 1160
-2.348777961004764e+01, // 1161
-4.714304332163732e+01, // 1162
 1.053573565902648e+01, // 1163
-1.107834996647511e+00, // 1164
 5.937321792714101e+01, // 1165
-3.667562829645500e+01, // 1166
 5.400749049767003e+01, // 1167
 1.283580161595815e+02, // 1168
-1.061210378760528e+01, // 1169
-7.629305449667213e+01, // 1170
 1.609088728336332e+01, // 1171
 1.801878628387392e+01, // 1172
-3.197036033265001e+01, // 1173
-1.053926289881935e+01, // 1174
-1.341587425188433e+01, // 1175
 3.126875061831739e+01, // 1176
-1.279566047506608e+01, // 1177
 9.891775302993116e+01, // 1178
-7.733470383674323e+00, // 1179
 8.079407972147559e+00, // 1180
 1.267671736672078e+01, // 1181
 2.497783188265934e+00, // 1182
 2.836321404487355e+01, // 1183
-4.063720993769122e+01, // 1184
-3.033148487625416e+01, // 1185
 4.797491769559025e+01, // 1186
-8.741189681895025e-01, // 1187
 1.303714896656780e+01, // 1188
-6.708883951781527e+01, // 1189
-3.335624632341597e+01, // 1190
 1.366266096360145e+01, // 1191
 3.055061316415479e+00, // 1192
 1.942338409192231e+01, // 1193
 1.384637787707477e+01, // 1194
-8.521201057431801e+01, // 1195
 1.201721161078134e+01, // 1196
-4.314297225998544e+01, // 1197
-2.583352444333000e+01, // 1198
 4.522996463793700e+01, // 1199
-4.063832718421800e+01, // 1200
-3.238857643339085e+01, // 1201
 2.964580661500252e+00, // 1202
 2.322141105352294e+01, // 1203
 2.975260488934033e+00, // 1204
-1.733405632618175e+01, // 1205
 2.298722443973154e+00, // 1206
-8.887897335761338e+00, // 1207
-1.652597395326459e+01, // 1208
 1.094540314162993e+02, // 1209
 5.824635870219440e+00, // 1210
-4.310785851610704e+00, // 1211
-1.124322074007168e+01, // 1212
-3.833346829813699e+00, // 1213
 2.967206251410087e-01, // 1214
 6.459657773894294e+00, // 1215
 6.736949611192424e+00, // 1216
-3.534016975887427e+01, // 1217
-1.051169339198311e+01, // 1218
-6.875998489334182e+00, // 1219
-1.221124183500750e+01, // 1220
-1.238686455670651e+01, // 1221
-1.266770642275900e+01, // 1222
 3.407118918826770e+00, // 1223
-9.277876606999362e+00, // 1224
-4.864718356176148e+00, // 1225
 8.631538502798783e+00, // 1226
-2.670963075017166e+00, // 1227
 8.850006055852166e+00, // 1228
 1.630624566732447e+01, // 1229
 6.052651712799441e+00, // 1230
 3.062784689831671e+01, // 1231
 5.763663153557515e+00, // 1232
-1.960997777452862e+01, // 1233
-1.590734231296642e+01, // 1234
 1.298592999477803e+01, // 1235
 3.242838878350194e+01, // 1236
 1.585792699505834e+01, // 1237
 7.456957187041716e+00, // 1238
-7.289938235280115e+01, // 1239
-2.116331337982208e+01, // 1240
-7.676031102505196e+01, // 1241
-4.173074591605767e+00, // 1242
 6.522676064652549e+01, // 1243
-5.011100073567444e+01, // 1244
 4.172549636018245e+01, // 1245
-1.634901479734393e+01, // 1246
-1.655506911032420e+00, // 1247
-3.397155590590918e+01, // 1248
-7.928155987512170e+01, // 1249
 3.509215954121236e+00, // 1250
-4.328033940798451e+01, // 1251
 3.094712502570069e+01, // 1252
-1.282069397795596e+02, // 1253
 1.706486348108102e+01, // 1254
 4.604336081247615e+01, // 1255
 5.049164173753283e+01, // 1256
 4.137032293569537e+01, // 1257
 1.032068089589036e+01, // 1258
 8.677948038754593e+01, // 1259
 4.568490520492595e+01, // 1260
-7.195962231807260e+01, // 1261
-9.122152652989338e+01, // 1262
-5.414997150198622e+01, // 1263
-3.341921486487182e+01, // 1264
-1.128394049554144e+01, // 1265
 2.059501669836411e+01, // 1266
-3.741530752524812e+01, // 1267
-3.123501059621393e+01, // 1268
-1.181821922532332e+01, // 1269
-3.380845567622274e+01, // 1270
 5.012924205079354e+01, // 1271
 7.122805587358050e+01, // 1272
-2.192035043159143e+00, // 1273
-2.676832162158393e+00, // 1274
 2.375430804465116e+01, // 1275
 5.194821246785191e+00, // 1276
-1.558188892729153e+01, // 1277
-2.290522253524860e+01, // 1278
-5.067344830848202e+00, // 1279
 1.378896906751466e+01, // 1280
 1.548759361816799e+01, // 1281
 5.393819465283518e+01, // 1282
-2.286879193450880e+00, // 1283
 1.820563599854976e+01, // 1284
 2.119704531052606e+01, // 1285
 4.738812555812678e+01, // 1286
-6.227873102563060e+00, // 1287
-3.914045299565406e+01, // 1288
 4.057001549659964e+01, // 1289
 3.427839243909359e+01, // 1290
-2.802492675406109e+01, // 1291
-3.294523677557743e+01, // 1292
 9.723598601441006e+00, // 1293
-1.067726346600404e+01, // 1294
-4.833396871816592e+01, // 1295
 7.019955157418622e+01, // 1296
-5.345808678748676e+01, // 1297
 6.917950559129442e+01, // 1298
 2.334476415988335e+01, // 1299
-3.295257265592478e+01, // 1300
-9.495663174998604e+01, // 1301
 4.544419034237494e+01, // 1302
-7.730612020633246e-01, // 1303
 3.203840602894491e+01, // 1304
 1.002359984962910e+02, // 1305
-2.553697492126233e+00, // 1306
-7.080897614212384e+01, // 1307
-1.466156258118231e+01, // 1308
 2.217497805853408e+02, // 1309
-7.788027428891472e+00, // 1310
-1.520283432037006e+02, // 1311
-3.062026439647300e+01, // 1312
-4.465033107772661e+01, // 1313
-5.563730844515288e+01, // 1314
-3.966936161000838e+01, // 1315
-1.747274101794914e+01, // 1316
-1.433454674320478e-01, // 1317
-6.319611609849379e+00, // 1318
 1.758788649660100e+01, // 1319
-3.805515238039199e+01, // 1320
-4.005266348442879e+01, // 1321
-7.323904474873508e+01, // 1322
-9.676999122449840e+01, // 1323
 1.001092310324462e+02, // 1324
-1.379957941682539e+01, // 1325
 1.548690871477634e+02, // 1326
 9.252525478787275e+01, // 1327
-6.524406895529290e+01, // 1328
 1.287044420546826e+01, // 1329
-3.678551946754342e+01, // 1330
 1.371568237668746e+00, // 1331
-1.999448602694672e+00, // 1332
 4.568910141471439e+00, // 1333
-1.435151202675838e+01, // 1334
 2.550318491279598e+01, // 1335
 5.762739589768380e+00, // 1336
-5.766299243937299e+01, // 1337
 7.655055118411351e+00, // 1338
-1.070247109003127e+02, // 1339
-2.981261350090351e+01, // 1340
-4.758708896539634e+01, // 1341
 9.992167276216043e+01, // 1342
 4.881179127569618e+00, // 1343
-1.570179003283429e+01, // 1344
 9.249580371096508e+01, // 1345
 8.058304415916852e+01, // 1346
-1.168674253566550e+02, // 1347
 4.510194131491696e+01, // 1348
-4.500627648414043e+01, // 1349
 2.381605206445117e+01, // 1350
-1.531099944639901e+01, // 1351
-3.999090400244751e+00, // 1352
 1.324263176375093e+02, // 1353
 1.014316322894901e+02, // 1354
 4.708749890410198e+01, // 1355
-1.879915542912514e+01, // 1356
-7.464870516997922e+01, // 1357
-1.714046084969060e+01, // 1358
-9.798537379100772e+01, // 1359
 1.645988911035696e-01, // 1360
-1.753891103672526e+01, // 1361
 4.648203583788645e-01, // 1362
 4.092570964341525e+01, // 1363
-2.583189495931681e+01, // 1364
-1.044845611251207e+00, // 1365
 4.218422088558049e+00, // 1366
-2.215169587126186e+01, // 1367
-2.163556955735882e+01, // 1368
-1.117716119588389e+01, // 1369
-2.080384465813374e+01, // 1370
-3.605240702140023e+01, // 1371
-1.359457442631426e+01, // 1372
-3.719843406151699e+00, // 1373
-9.480399590721223e+00, // 1374
-2.202637495107123e+00, // 1375
-1.133410659292543e+00, // 1376
 3.484751487246013e+01, // 1377
 3.253505686617715e-01, // 1378
 5.149661369829450e+00, // 1379
 3.976766011141367e-01, // 1380
-3.892312965077107e+01, // 1381
-8.889632798345417e+00, // 1382
-1.620006260366527e+01, // 1383
-1.997625528088289e+00, // 1384
-4.483239406668226e+00, // 1385
-1.732801111067309e+00, // 1386
-7.883904027548749e+00, // 1387
-2.954649818498381e+01, // 1388
-4.052820804430097e+00, // 1389
-4.381969587312386e+00, // 1390
-2.953971117128739e+00, // 1391
-8.729940216507406e-01, // 1392
 1.201851191897509e+00, // 1393
 7.528696978593627e+00, // 1394
 1.877075449085862e+00, // 1395
-2.811912287917756e+01, // 1396
-6.204806140006530e+00, // 1397
-1.978918789920972e+01, // 1398
-5.559806243486109e+00, // 1399
-7.146757230252969e+00, // 1400
-3.904278951232158e+00, // 1401
-1.646345801014036e+00, // 1402
-4.931949566487615e+00, // 1403
 4.958210266517870e+01, // 1404
-1.778349834617232e+01, // 1405
-3.563120665777689e+01, // 1406
-1.638369377060750e+01, // 1407
-2.023627426600692e-01, // 1408
-2.684811297669885e-01, // 1409
-1.244591214834695e+00, // 1410
-4.322773221032193e-01, // 1411
 1.204548583406671e+00, // 1412
-1.471744117963699e+00, // 1413
-5.621848404717873e+00, // 1414
-1.115625707080266e+00, // 1415
-1.274237982614864e+01, // 1416
-3.570210563443207e+01, // 1417
-5.541488756114885e+00, // 1418
-4.208229385171152e+00, // 1419
-3.802621908078060e+00, // 1420
-3.187885688163051e+00, // 1421
 1.289373937868621e+00, // 1422
 4.678849141933230e+00, // 1423
 1.640111609421334e+00, // 1424
-3.085182433040482e+01, // 1425
-6.341343923962429e+00, // 1426
-2.479330547470478e+01, // 1427
-6.181850507433975e+00, // 1428
-8.437679227284477e+00, // 1429
-8.976380796076512e+00, // 1430
-2.553394792753108e+00, // 1431
-6.790915658024709e+00, // 1432
-4.063071907244571e+01, // 1433
-5.943217737121634e-01, // 1434
-2.872636099223288e+01, // 1435
-4.808933169175898e-01, // 1436
-5.239240601885600e+00, // 1437
-4.339788711723582e+00, // 1438
-1.906369400213591e+00, // 1439
-8.485130501638526e+00, // 1440
 2.228111970153167e+01, // 1441
-9.785686067786109e+01, // 1442
 3.214805340080405e+01, // 1443
-2.723781046868998e+01, // 1444
-9.906603306758790e+01, // 1445
 7.500818092462913e+01, // 1446
-4.890900131271024e+01, // 1447
 8.529949830575848e+01, // 1448
 5.109600624213165e+01, // 1449
 7.171695481145151e+00, // 1450
-4.443585055462106e+01, // 1451
-8.623886872500714e+00, // 1452
 1.081746995496791e+02, // 1453
-1.621963316363802e+01, // 1454
-2.203859368571679e+01, // 1455
 3.015224453416431e+01, // 1456
 7.420158176666553e+01, // 1457
-3.054430424469784e+01, // 1458
-1.204257959583021e+02, // 1459
 3.221090980247038e+01, // 1460
-1.749957061654329e+01, // 1461
-5.217390501174870e+01, // 1462
-1.188784308955628e+02, // 1463
 9.147664097429389e+01, // 1464
 3.162120826959145e+01, // 1465
 7.167467797448911e+01, // 1466
-1.766290658788190e+01, // 1467
 1.678480359430059e+02, // 1468
 4.047406873948385e+01, // 1469
 8.872874934674625e+00, // 1470
-8.326902253123082e+01, // 1471
 6.202066967583178e+01, // 1472
 2.215157786167340e+02, // 1473
 1.517277949857418e+02, // 1474
 1.981501802470445e+02, // 1475
 3.027294117003465e+00, // 1476
-1.653147557706807e+02, // 1477
-3.468612146951953e+01, // 1478
 2.292009882316454e+01, // 1479
-2.282643890056480e+01, // 1480
 6.817070374523358e+01, // 1481
-1.251025972406577e+02, // 1482
 2.497084788062795e+02, // 1483
 1.969824742932965e+02, // 1484
 8.946775360351629e+01, // 1485
-1.407542811892008e+02, // 1486
-3.728870153854958e+01, // 1487
-2.126259057078967e+00, // 1488
-9.244025604029228e+01, // 1489
 6.530296344379021e+00, // 1490
 1.303404124609293e+01, // 1491
-8.864256291105276e+01, // 1492
 1.239500440382744e+02, // 1493
 2.383281991299824e+01, // 1494
 1.323705740296197e+02, // 1495
-1.467025803486329e+00, // 1496
-5.353993171144266e+01, // 1497
 1.483723028248731e+02, // 1498
-6.765158090374952e+01, // 1499
 8.358574874431180e+01, // 1500
 1.859706356923026e+01, // 1501
 2.927128186210815e+01, // 1502
-4.835021132800267e+01, // 1503
 4.191669594322022e+01, // 1504
-1.134710715870091e+02, // 1505
-6.640640856176777e-01, // 1506
 8.199030633303221e+01, // 1507
-3.631671447573331e+01, // 1508
-1.989961359868975e-03, // 1509
-3.310534170434514e+01, // 1510
-1.225057879176537e+01, // 1511
 3.717446140345900e+01, // 1512
 6.983376988806474e+01, // 1513
 1.589083377271470e+01, // 1514
 9.851629041207850e+00, // 1515
 1.039138640569047e+01, // 1516
-6.087278172651109e+01, // 1517
-3.096920563135616e+01, // 1518
 3.902078833284622e+01, // 1519
-9.986324059562855e+01, // 1520
 3.613835731348183e+01, // 1521
-1.197447364870659e+01, // 1522
 3.603215246529716e+01, // 1523
-1.718896750750770e+02, // 1524
 5.522331967318799e+01, // 1525
-4.232899838605183e+00, // 1526
 1.027428356669293e+02, // 1527
-8.151497104724736e+01, // 1528
-3.921884671248916e+01, // 1529
-7.377727894923902e+01, // 1530
 4.913453118752394e+01, // 1531
 9.813773133870407e+01, // 1532
 9.618900483990802e+01, // 1533
 1.984637570914872e+01, // 1534
 8.706201181768254e+00, // 1535
-9.689933029177899e+01, // 1536
 6.721207692546223e+01, // 1537
 3.313211650923017e+01, // 1538
 7.954544420712975e+01, // 1539
 5.815137435433240e+01, // 1540
 1.272820854040791e+02, // 1541
 7.761925939746322e+01, // 1542
 4.319424866373491e+01, // 1543
 4.447176258801917e+01, // 1544
-4.544083202363145e+01, // 1545
-5.190700496769128e+01, // 1546
 1.461800413627847e+01, // 1547
-5.384080108629470e+01, // 1548
-1.521527509941720e+01, // 1549
-2.617560019768083e+01, // 1550
-1.382974292585761e+02, // 1551
-1.479433079173150e+02, // 1552
 6.990886283859651e+01, // 1553
 7.787633098130708e+01, // 1554
 4.534164570406798e+01, // 1555
-1.624741733247642e+02, // 1556
-1.431606262518989e+01, // 1557
-1.556650504071544e+02, // 1558
-4.495501545515111e+01, // 1559
-2.926410134499866e+01, // 1560
 3.438855138435697e+01, // 1561
 6.153953407969473e+01, // 1562
-6.433912028044777e+01, // 1563
 1.244447107018692e+01, // 1564
-2.235994033382350e+01, // 1565
 1.472341151677923e+01, // 1566
 8.550464502030394e+01, // 1567
-7.217245825296996e+01, // 1568
-7.165688534980373e+00, // 1569
 9.376023979366673e+00, // 1570
-7.973439001242396e+01, // 1571
-2.451935336028632e+01, // 1572
 1.910414141990627e+01, // 1573
-9.582949844794010e+01, // 1574
-2.062513889819948e+00, // 1575
-2.874282329758691e+01, // 1576
 7.478528201186464e+01, // 1577
 4.675357127729725e+01, // 1578
 7.232937983504016e+00, // 1579
-1.126126312627703e+02, // 1580
 2.349029561235534e+01, // 1581
-2.786047294122097e+01, // 1582
-3.687169128441734e+01, // 1583
 1.259087119270662e+01, // 1584
 2.166978737108753e+01, // 1585
 7.210906571250135e+01, // 1586
-2.146988947172199e+02, // 1587
-5.598025854253554e+00, // 1588
-4.942079670023015e+01, // 1589
-2.590145868813638e+01, // 1590
 6.301988655011352e+01, // 1591
 1.572047969833938e+01, // 1592
-1.054501248859052e+02, // 1593
 4.510475788966259e+01, // 1594
-1.452312014443856e+01, // 1595
 5.294154023325151e+00, // 1596
 1.093795426707236e+02, // 1597
 4.631995899891755e+01, // 1598
 1.076270689511039e+01, // 1599
-4.686961242149766e+01, // 1600
-6.174786898160446e+01, // 1601
 2.912006024181414e+01, // 1602
-3.924948393685782e+00, // 1603
 4.964180099921804e+01, // 1604
-9.155502933226650e+00, // 1605
 4.110092413259120e+01, // 1606
-4.548543202930514e+00, // 1607
-1.698448975849939e+02, // 1608
 6.833955430942656e+01, // 1609
-7.899522373372233e+01, // 1610
 2.843332375682661e+01, // 1611
-3.381220393285512e+00, // 1612
 4.535394697871865e+00, // 1613
-2.198198310272368e+02, // 1614
-1.383650814165851e+01, // 1615
 3.229197469047229e+00, // 1616
-2.518617469172522e+02, // 1617
-3.015376395245806e+01, // 1618
-2.080392960758211e+01, // 1619
 2.193672453363321e+01, // 1620
 2.504893314130531e+01, // 1621
-1.124370880163414e+02, // 1622
 4.170058181571212e+01, // 1623
-1.344283738855945e+00, // 1624
-2.900364071358859e+00, // 1625
-2.306106082743910e+01, // 1626
-1.352118861815050e+01, // 1627
-3.919015801231834e+01, // 1628
 1.668699898644756e+01, // 1629
-1.073967024596228e+02, // 1630
 1.063272592034703e+02, // 1631
 2.430901887466717e+00, // 1632
-1.347631335179141e+01, // 1633
 5.050629073321830e+01, // 1634
 9.962291916480440e+00, // 1635
-4.437054885070666e+01, // 1636
 5.292324420144272e+01, // 1637
 5.481897364608280e+01, // 1638
-3.102581907325830e+01, // 1639
-4.952152405063136e+00, // 1640
-5.423470464040052e+01, // 1641
 4.594994065241915e+01, // 1642
 7.381197804573709e+01, // 1643
 7.718220760696147e+00, // 1644
-1.986352063946448e+01, // 1645
 4.351018677174666e+01, // 1646
 1.870983528259745e+02, // 1647
 1.165406457609850e+02, // 1648
-1.057969799576449e+01, // 1649
 3.180075817627018e+02, // 1650
 5.725335536694935e+01, // 1651
-1.705169425943444e+01, // 1652
-1.376427079718897e+02, // 1653
-3.315749107030546e+01, // 1654
 4.590945121902364e+01, // 1655
-5.312544878785862e+01, // 1656
 3.091811519017369e+01, // 1657
-9.798316947442281e+01, // 1658
 3.936220032699736e+00, // 1659
 7.062686703990714e+01, // 1660
 2.798663783214814e+01, // 1661
 1.101797932635545e+02, // 1662
-9.101768286671805e+01, // 1663
 3.132410423376215e+01, // 1664
-8.104626588450999e+01, // 1665
-7.998699607576816e+01, // 1666
-8.390023294526517e-01, // 1667
 6.550158849089224e+00; // 1668

}

netcdf mbnrg_2b_A1B3C1D2_E1F2_fit {
  // global attributes 
  :name = " mbnrg_2b_A1B3C1D2_E1F2_fit";
  :k_x_intra_A_B_1 =  3.313005746029803e-01; // A^(-1))
  :k_x_intra_A_C_1 =  4.401841146487998e-01; // A^(-1))
  :k_x_intra_A_D_1 =  2.461155200940438e+00; // A^(-1))
  :k_x_inter_A_E_0 =  8.571191506394328e-01; // A^(-1))
  :k_x_inter_A_F_0 =  2.261519988786035e-01; // A^(-1))
  :k_x_intra_B_B_1 =  1.849899959001211e+00; // A^(-1))
  :k_x_intra_B_C_1 =  1.880179488341646e+00; // A^(-1))
  :k_x_intra_B_D_1 =  2.632342848980163e-01; // A^(-1))
  :k_x_inter_B_E_0 =  7.739478000384370e-01; // A^(-1))
  :k_x_inter_B_F_0 =  6.912877955728575e-01; // A^(-1))
  :k_x_intra_C_D_1 =  5.812702756358955e+00; // A^(-1))
  :k_x_inter_C_E_0 =  1.180195341744499e+00; // A^(-1))
  :k_x_inter_C_F_0 =  9.457780848959891e-01; // A^(-1))
  :k_x_intra_D_D_1 =  2.393509279645449e+00; // A^(-1))
  :k_x_inter_D_E_0 =  4.812296137910029e+00; // A^(-1))
  :k_x_inter_D_F_0 =  6.000375011983535e-01; // A^(-1))
  :k_x_intra_E_F_1 =  4.195649209887358e-01; // A^(-1))
  :k_x_intra_F_F_1 =  2.599849643205974e+00; // A^(-1))
  :ri =  6.000000000000000e+00; // A
  :ro =  7.000000000000000e+00; // A
  dimensions:
  poly = 1183;
  variables:
    double poly(poly);
data:
poly =
 7.868784220337318e+01, // 0
 1.271106915227615e+02, // 1
-2.171405714768526e+02, // 2
 1.075063077255816e+02, // 3
 2.146888122182886e+01, // 4
-1.263013432921046e+02, // 5
-2.799235879241697e+02, // 6
 2.876228147575003e+01, // 7
 1.633893440486446e+02, // 8
 3.001638832562597e+02, // 9
-1.005218066300646e+00, // 10
-3.148311341478610e+02, // 11
-2.820888760510354e+02, // 12
 2.119508602278733e+02, // 13
 3.685747956119222e+01, // 14
 2.192820199000511e+02, // 15
 1.555104422048608e+02, // 16
-7.936876693076168e+01, // 17
-1.409154014110283e+02, // 18
-1.212198243962192e+02, // 19
-1.440560151016507e+01, // 20
 2.683240846875800e+02, // 21
 1.203960284400854e+02, // 22
 4.248020000169585e+02, // 23
 5.534734887666944e+00, // 24
 5.412042892217778e+02, // 25
 2.782032868119621e+02, // 26
 3.999722920160623e+00, // 27
 1.785941448208297e+02, // 28
 1.769801264130978e+02, // 29
 4.827396834680698e+01, // 30
 9.442834578239899e+01, // 31
 3.096183392147264e-01, // 32
 4.753028423456238e-03, // 33
 3.970312075735754e-01, // 34
 2.708537163586067e+02, // 35
 1.904399579346601e+00, // 36
 1.754895747866658e+02, // 37
 1.713571732419414e+02, // 38
 9.291246297307484e+01, // 39
 9.079954174638597e+01, // 40
 4.235623397237367e-01, // 41
 3.047702348217197e+01, // 42
 1.035180991995098e+02, // 43
-2.002290999429458e-01, // 44
-9.878069036154112e-03, // 45
-2.481836039831417e-01, // 46
 8.222946770554915e-02, // 47
 9.716642310138156e-04, // 48
-2.305570811181235e-01, // 49
-1.732117200914910e-03, // 50
 7.193133100545964e+01, // 51
-3.431170060677346e+02, // 52
-3.807497776710702e+02, // 53
 1.187953198790751e+02, // 54
 2.323090103558249e+02, // 55
-5.293208431567352e+00, // 56
-1.677401156946788e+00, // 57
 4.579657864491383e-03, // 58
-3.052447353785740e+00, // 59
-3.937959189889300e-02, // 60
 2.784322701533623e+02, // 61
-2.006437019812417e+02, // 62
 1.879441799494715e+02, // 63
-2.962439951907190e+02, // 64
 7.334177847874365e+01, // 65
-2.712321564440723e+02, // 66
 1.224170675161293e+02, // 67
-7.425551292008962e+02, // 68
-3.854511213974507e+02, // 69
-3.345682662646057e+02, // 70
-1.555569131575061e+02, // 71
 1.587235744124926e+02, // 72
-7.260753602039794e+01, // 73
 7.025213628029801e+02, // 74
-2.226708704363033e+02, // 75
-3.480527697941494e+02, // 76
-6.702403330678833e+02, // 77
 1.061079107246881e+03, // 78
 9.225426850524003e+01, // 79
 1.019124119186096e+00, // 80
 6.065976982019266e+01, // 81
 5.814705039252096e+01, // 82
 4.078700157730468e+01, // 83
 3.505500797080852e+01, // 84
 8.152275409161407e-02, // 85
 2.789616585028337e+01, // 86
 3.285156242018911e+01, // 87
-7.760869641170524e-02, // 88
 4.157617246391187e+01, // 89
 7.094763173213458e+01, // 90
-4.292056829505960e+01, // 91
-1.116339861655463e+00, // 92
-1.332783651036938e+01, // 93
-2.431174744653953e+01, // 94
-1.004220768669197e+02, // 95
-1.803855857671168e+02, // 96
 8.307044311791470e+00, // 97
 1.133977433725328e+01, // 98
-3.601534884474804e+02, // 99
 1.151918453057392e+02, // 100
-1.495776897789220e+02, // 101
 8.170534953832812e+02, // 102
 7.628924305096417e+02, // 103
 3.004209601274459e+02, // 104
 1.140794390565272e+01, // 105
 8.797365945644960e+01, // 106
 4.661909667753682e+02, // 107
 2.715247806182667e+02, // 108
-2.936743529455489e+02, // 109
 9.373626194285978e+01, // 110
-3.825738946301814e+01, // 111
-2.552065416865163e+02, // 112
-1.717557407815446e+01, // 113
-1.311557103119351e+02, // 114
-5.221854831416454e+02, // 115
 8.428039117790921e+02, // 116
 4.822169163576928e+02, // 117
-2.875879433803233e+02, // 118
 2.095247094471086e+02, // 119
 7.322255707452200e+01, // 120
 1.154413105161149e+00, // 121
 9.465841652676217e+01, // 122
 4.519098713454433e+01, // 123
 4.459614867703999e-02, // 124
 4.577251790519641e+01, // 125
 3.068384801454279e-02, // 126
-5.820214673391015e+01, // 127
-1.604660962020662e+02, // 128
 8.095165230024451e-03, // 129
-4.885276414218189e+01, // 130
 8.259525261867287e+00, // 131
 7.384752964052277e+01, // 132
-1.671663667202460e+02, // 133
 3.917712798373779e+02, // 134
-1.872048311465587e+02, // 135
 1.711754271590907e+01, // 136
 4.032832496473524e+00, // 137
 2.431759237082474e+02, // 138
 2.593017732759695e+02, // 139
 2.793648341490776e+02, // 140
 5.600012768033677e+00, // 141
 3.432364270959185e+02, // 142
 1.339844483301523e+03, // 143
 1.163808955541784e+01, // 144
-4.376522022368594e+01, // 145
 3.461974851058247e+02, // 146
 3.526634651127708e+02, // 147
 1.342794718103879e+02, // 148
 2.639811482266729e+01, // 149
-4.395945133213514e+01, // 150
 5.653908239733166e-01, // 151
 2.589505958143423e-01, // 152
-1.991566247720905e-03, // 153
-1.368816122896263e+02, // 154
-1.284613288727288e+02, // 155
-1.414896436033124e+02, // 156
 3.176177434475532e-01, // 157
-4.521516677360282e+01, // 158
-2.784618006419123e+01, // 159
-7.563677411607350e-01, // 160
-7.544189999364843e-02, // 161
 1.089296240358105e-03, // 162
-1.983000098999960e-01, // 163
-2.527223662866429e-03, // 164
-1.183166117348572e+02, // 165
-2.095818578682791e+01, // 166
-9.695551191709511e+01, // 167
 1.160163938666144e-01, // 168
-4.982571569665232e+01, // 169
-7.385718170500343e+01, // 170
-8.906983473721314e-02, // 171
-1.194847735116094e+01, // 172
-8.321770481108001e+01, // 173
 1.436754893174313e+02, // 174
 1.286016333754619e+01, // 175
 1.329718197714331e-01, // 176
-3.264528321419091e+01, // 177
-1.998160062451939e-02, // 178
-1.204721952754172e+00, // 179
-7.776902473868398e-01, // 180
 2.351175345206164e+01, // 181
 1.566794472118484e+02, // 182
-1.042391732161535e+02, // 183
 7.911211161402935e+01, // 184
 1.924461378837520e+02, // 185
-2.652611104529831e+02, // 186
-4.232321535328219e+01, // 187
-4.328671538245802e+02, // 188
 3.503139637590439e+02, // 189
 3.223801187399427e+01, // 190
-3.587150975325713e+02, // 191
-1.435844670818749e+02, // 192
-6.450876083700194e+01, // 193
 1.297820749793258e+02, // 194
-2.941786545155934e+01, // 195
-2.317459501142324e+02, // 196
-2.279272253329225e+02, // 197
-6.476113232628067e+01, // 198
 1.518086249822081e+02, // 199
-5.421058361846754e-01, // 200
 9.578108763251684e+01, // 201
 9.915405890931699e+01, // 202
 8.265101041424099e+01, // 203
 6.126353420664206e+01, // 204
 1.337746890704776e-01, // 205
 5.474963669874446e+01, // 206
 4.323157092058024e+01, // 207
-4.630868549487280e-01, // 208
 2.451343009842455e+01, // 209
 1.570160422383816e+02, // 210
 7.596608279489300e+01, // 211
-8.528861282975141e+00, // 212
-1.862425903595233e+00, // 213
 1.556040431015606e+01, // 214
 1.340738226508484e+01, // 215
-1.878277722438323e+02, // 216
 2.329345680327053e+01, // 217
 2.309851125738219e+02, // 218
 3.503985503171153e+01, // 219
 1.143009587546861e+02, // 220
 8.021133691706018e+01, // 221
-2.369934871172865e+02, // 222
 6.204781001980973e+00, // 223
 3.145374815586318e+01, // 224
 6.290781178966574e+02, // 225
-5.625172308884230e+02, // 226
 3.586882365649557e+02, // 227
 1.229890988543081e+01, // 228
 2.890427064623281e+02, // 229
 1.437038575409269e+02, // 230
-2.433167233044227e+02, // 231
 2.686680165609681e+02, // 232
-7.545097854127850e+01, // 233
 2.373390647214015e+01, // 234
 1.794529795303020e+02, // 235
 5.236870592940777e+02, // 236
-6.253712132363322e+02, // 237
 3.155816704147140e+01, // 238
 1.253935015578720e+02, // 239
 6.076072475692322e+02, // 240
 7.872914997983199e+01, // 241
 4.367945569686242e+02, // 242
 2.432334324008720e+01, // 243
 7.797419776966076e+01, // 244
 7.974818584771319e+00, // 245
 7.038065691974349e-03, // 246
 1.464451033072684e+02, // 247
 1.298183252671920e+02, // 248
-8.472766442551792e-01, // 249
 5.475156561042653e+01, // 250
 3.627182417253391e+00, // 251
 9.444857112677502e+01, // 252
-3.376302359947467e+01, // 253
 3.598798834546086e+01, // 254
 1.291931267647952e+02, // 255
-2.998396908084920e+01, // 256
 1.259770481269213e+01, // 257
 1.886705995810421e+02, // 258
-9.191011258195007e+01, // 259
-9.805084331168587e+00, // 260
-4.794066834881602e+01, // 261
-2.524579280638799e+02, // 262
 1.037751775863341e+01, // 263
-7.135234258379337e+01, // 264
-6.575135086177147e+01, // 265
 9.979415560582386e+01, // 266
-2.909599397995444e+02, // 267
 1.147599595415591e+01, // 268
-2.177363720935255e+02, // 269
 6.432852804182082e+01, // 270
-4.611281194801953e+01, // 271
 2.734537594287521e+02, // 272
-7.419100868739211e+01, // 273
 7.992606096598396e+01, // 274
 5.120031349839740e+02, // 275
-1.331496850400531e+01, // 276
 1.038263135160488e+01, // 277
 7.738652821031275e+01, // 278
-6.745545057644402e+01, // 279
 8.942963835712288e+00, // 280
 1.000090816409092e+02, // 281
 1.009558172581513e+02, // 282
-4.464570358249268e+02, // 283
-1.179047193899649e+01, // 284
-1.751233147972364e+02, // 285
-1.503894456302539e+01, // 286
 3.175988875548856e+01, // 287
 1.190096139274112e+02, // 288
 3.431391062084685e+02, // 289
 2.048731742705919e+02, // 290
 2.903520316481962e+01, // 291
 1.905040825352906e+01, // 292
-1.275300980741715e+02, // 293
 2.268133369892427e+02, // 294
-5.997413889652842e+01, // 295
-4.503212882710338e+02, // 296
-4.490759811784148e+00, // 297
-1.178725252533372e+02, // 298
 4.090345597625359e+02, // 299
-2.353616455847538e+02, // 300
 7.481008440381584e+02, // 301
-5.020086912948495e+01, // 302
-6.962519144044560e+01, // 303
 1.180890687568452e+01, // 304
 3.739679106925271e+02, // 305
 3.909141176649676e+02, // 306
 1.086301034600428e+01, // 307
 8.173650491577656e+01, // 308
 1.594125255905352e+02, // 309
-2.632384316132693e+02, // 310
-1.490582841415648e+02, // 311
 1.641514040988454e+02, // 312
 1.281371717941160e+02, // 313
 1.386462193952886e+00, // 314
 1.652409446745108e+02, // 315
 7.442549634062897e+01, // 316
 6.762328210625365e-02, // 317
 7.942477003789843e+01, // 318
-4.972822562117613e-02, // 319
-7.758416786808178e+00, // 320
-5.268188500201324e+01, // 321
-2.716304596259799e+00, // 322
-6.106232036121989e+00, // 323
 2.446718907092006e+02, // 324
 3.132517865263112e+02, // 325
-4.513663591741704e+02, // 326
 1.522607929423744e+01, // 327
-3.701971118142585e+02, // 328
 3.189984079685798e+01, // 329
 2.807516041253132e+02, // 330
 8.311349424431951e+01, // 331
-3.648903793318568e+02, // 332
 1.097459032022481e+02, // 333
 7.759882071232468e+01, // 334
-1.675578362224603e+02, // 335
 9.375290181376045e+02, // 336
 2.229667603608128e+01, // 337
 1.874342850844249e+01, // 338
 7.175996418787325e+01, // 339
 2.997670560167960e+02, // 340
 2.072864342692986e+02, // 341
 3.331023788317501e+01, // 342
-5.378519245921584e-02, // 343
 1.168540128368686e+02, // 344
-2.365320173676838e-01, // 345
 8.408008921258009e+01, // 346
 3.717282342523909e+01, // 347
 9.348563052464914e+01, // 348
-2.468478574414778e+02, // 349
 2.377728657600217e+02, // 350
-2.672457471318920e+02, // 351
 2.077566002887547e+02, // 352
-1.330447864177586e+02, // 353
 4.104445365494063e+01, // 354
-1.333719329812025e+02, // 355
-4.440435125525335e+01, // 356
 4.122654917713488e+02, // 357
 1.754352418029995e+02, // 358
-1.364215201088402e+02, // 359
 9.242414989430907e+01, // 360
 3.367309865710033e+02, // 361
-2.426605527307514e+01, // 362
-2.710626869448411e+02, // 363
-3.979015416177755e+01, // 364
 1.675337300824048e+01, // 365
 3.106035545362242e+02, // 366
-1.504643589133914e+02, // 367
 1.117559626544632e+01, // 368
-3.258267115552726e+01, // 369
 2.292587658268483e+02, // 370
 1.099455766850427e+02, // 371
-5.323945984261866e+01, // 372
-5.825559878758784e+02, // 373
-2.812447984465244e+02, // 374
-3.313787144504792e+01, // 375
 1.172851475194693e+02, // 376
-4.454598725917658e+02, // 377
-3.830028589736680e+02, // 378
-4.487542005086133e+02, // 379
 2.404073122217253e+02, // 380
 2.753591380378266e+01, // 381
 2.841517055276008e+02, // 382
-1.204996866706175e+02, // 383
 3.515537156731783e+02, // 384
-7.570763826820812e+02, // 385
-4.192417828976427e+01, // 386
 7.387438744297920e+02, // 387
-4.927056919809709e+02, // 388
-1.812258467764136e+02, // 389
-6.088069147717346e+02, // 390
 3.373089510134653e+02, // 391
-1.119474590930970e+02, // 392
 1.152451162857716e+02, // 393
 3.180277143393197e+02, // 394
-2.529019250072689e+02, // 395
 1.465353268119664e+01, // 396
 1.682450719091488e+02, // 397
 4.106309070789208e+02, // 398
-3.278120724185931e+02, // 399
-5.981765969649248e+01, // 400
 1.575101884733675e+02, // 401
 9.396094255536741e+01, // 402
-5.455457269514095e+01, // 403
 6.513507423425551e+02, // 404
 3.522688442377471e+01, // 405
 1.986299348982121e+02, // 406
 3.078944757475609e+01, // 407
 6.641739272899617e+02, // 408
 4.265188430076646e+02, // 409
-2.918608737746540e-01, // 410
 5.896535379741011e+00, // 411
 1.509812590658804e+01, // 412
-3.297711483757578e+01, // 413
 4.087462548418538e+02, // 414
-3.159556666289572e+02, // 415
 1.725699272543320e+02, // 416
 6.931386809754442e+02, // 417
 4.440561958543806e+02, // 418
 8.948374492413783e-01, // 419
 4.410616790412543e+02, // 420
-3.235048519856414e-01, // 421
 5.961019956843929e+01, // 422
-3.025917693494042e-01, // 423
-1.078701140619351e+02, // 424
 1.427533552288221e+02, // 425
 3.779805492010273e+02, // 426
-5.438960405005976e+02, // 427
 1.570301959100156e+02, // 428
 6.943349994450182e+01, // 429
 1.538056149592532e+02, // 430
-1.107274981652732e+02, // 431
-4.341001481938138e+02, // 432
 1.123054462971469e+02, // 433
 4.494185309272571e+02, // 434
 1.149419444568487e+02, // 435
 7.665562828515480e+01, // 436
 6.483951234739054e+02, // 437
-2.170838446282586e+01, // 438
 2.376399876051588e+02, // 439
 2.573597137941311e+02, // 440
 1.800301635404611e+02, // 441
-1.535467426774910e+02, // 442
-3.121224590268582e+02, // 443
 1.530794568204282e+02, // 444
-1.385439509642555e+02, // 445
-1.871994137289510e+02, // 446
 1.380867998831188e+02, // 447
-9.470324683334870e+01, // 448
 1.877057379022668e+02, // 449
 9.293472552965835e+01, // 450
 5.026074502602770e+00, // 451
 8.368502170723220e+01, // 452
-3.922481205817188e+02, // 453
 1.335740596687584e+02, // 454
 5.868202876274174e+02, // 455
 1.243578823148609e+02, // 456
 1.883246166186852e+02, // 457
-1.606535323508153e+02, // 458
-1.236891322304426e+02, // 459
 1.381916362340003e+02, // 460
-1.347577814165700e+01, // 461
-1.530854340530417e+02, // 462
 1.331035583042804e+02, // 463
-4.220730745614707e+02, // 464
-2.171095652125360e+02, // 465
 8.716074614223767e+01, // 466
 3.828361526330567e+02, // 467
 4.703130701566414e+02, // 468
 7.763623056886124e+01, // 469
 2.992835071300611e+02, // 470
 3.533902922250808e+02, // 471
-1.029647442252476e+02, // 472
 2.666804894686263e+00, // 473
-8.700934764927965e+01, // 474
-5.690885886706535e+01, // 475
-2.715983341432758e+02, // 476
-1.184065011861267e+02, // 477
-1.316075258034477e+02, // 478
 5.686883481421032e+02, // 479
 6.516159511753132e+01, // 480
-1.041658456787413e+03, // 481
 6.390625404897197e+01, // 482
 1.623140930913458e+02, // 483
-2.718885531220906e+02, // 484
 2.393076388447735e+02, // 485
 7.593702510592721e+01, // 486
 3.522403869370788e+02, // 487
 7.301757623782184e+01, // 488
-7.212382531794756e+01, // 489
-2.201759503505047e+02, // 490
 1.188584518307613e+00, // 491
 8.585428071635566e+01, // 492
 2.564370605178999e+01, // 493
 2.273125544682270e+01, // 494
 1.507176250943609e+01, // 495
 1.589278438689650e-02, // 496
 1.611816700318362e+01, // 497
-2.044912708338658e-02, // 498
-2.391054566834517e+02, // 499
-8.210161055372453e+01, // 500
 2.634695186871818e+02, // 501
 5.420157108731565e+00, // 502
 4.322574890560383e+00, // 503
 1.881296701991314e+02, // 504
 8.442398529088236e+01, // 505
 6.719062951064650e+01, // 506
 4.039592780914480e+00, // 507
 3.920187928733837e+01, // 508
 2.909185040871888e+01, // 509
 1.116077991714857e+02, // 510
 6.146355409758148e+01, // 511
-1.266832684167807e+02, // 512
 5.936391694498064e+00, // 513
 1.743187834284569e+01, // 514
-9.450035432971500e+00, // 515
-3.692427592211776e+00, // 516
-4.366912389640004e+01, // 517
 1.344228379977475e+02, // 518
-1.980772985823756e+02, // 519
-2.020696377090038e+02, // 520
-4.263798898795248e+01, // 521
-1.476273001699487e+02, // 522
 3.716540310002288e+00, // 523
-2.946358021460365e+01, // 524
 8.246134563761750e+00, // 525
-4.984098679992454e+00, // 526
-1.381994007191846e+01, // 527
-3.142107707081240e+02, // 528
-3.358590907879793e+00, // 529
-6.394200299531758e+01, // 530
-4.705669853129744e+01, // 531
 2.312917833939140e+02, // 532
 2.091756397556264e+00, // 533
-1.656816999470655e+02, // 534
-7.835491180053214e+01, // 535
-2.131705451100382e+02, // 536
-4.708325916753998e+00, // 537
 4.986326406004967e+01, // 538
 1.452246896305866e+02, // 539
-5.407373546140808e+01, // 540
-1.768424611242897e+02, // 541
 9.243972616090561e+01, // 542
-4.021425239550903e+02, // 543
 1.522983818082945e+00, // 544
-2.524983416579720e+02, // 545
-1.575224196867820e+02, // 546
 4.585087316129059e+02, // 547
 2.614155921132186e+02, // 548
 3.756831156473445e+01, // 549
 1.521791227748317e+02, // 550
-1.437497181745823e+01, // 551
 1.169356244404382e+01, // 552
-1.462244704418615e+02, // 553
 4.884276884307681e+02, // 554
-8.504827238301360e+00, // 555
 6.399444263134691e+01, // 556
 3.220236793215062e+01, // 557
 3.059950574717701e-02, // 558
 3.721541681069071e+01, // 559
-2.470102520598182e-02, // 560
 2.499123214029862e+01, // 561
-6.042515305225005e+01, // 562
 5.833112720908164e+01, // 563
 9.428047620309613e+00, // 564
-5.866866483386302e+01, // 565
 4.271942643885217e+01, // 566
-3.286533394040685e+02, // 567
-3.672782490368402e+02, // 568
 8.837923965065078e+00, // 569
-3.054220222044693e+02, // 570
-3.536370820164591e+01, // 571
 1.095004115210259e+02, // 572
-3.372441508358341e+02, // 573
 1.831648453568063e+02, // 574
 4.210941023332322e+00, // 575
 4.517958282833512e+01, // 576
 3.771823723300020e+02, // 577
-2.314011187145774e+02, // 578
-1.109779422896278e+02, // 579
 4.476823447969977e+02, // 580
 1.089762610342136e+02, // 581
-4.018435674441908e+01, // 582
 4.839294425962064e+00, // 583
 4.061378109816856e+01, // 584
-5.186056310282510e+01, // 585
-3.881719604990306e+02, // 586
-3.376906637912210e+02, // 587
 4.073173839855200e+01, // 588
-3.745622952186648e+02, // 589
 2.460499865060675e+02, // 590
 1.232000752559751e+01, // 591
 3.689161825211392e+01, // 592
 2.600463161329626e+02, // 593
 4.342137770099632e+02, // 594
-3.473740069572215e+02, // 595
-2.608957072439899e+02, // 596
-2.288433996653367e+02, // 597
-1.483752833284955e+02, // 598
 3.028574024028349e+02, // 599
 2.351415700480090e+01, // 600
-1.578578622780939e+02, // 601
-3.144493197832211e+02, // 602
 2.188189944526532e+02, // 603
 1.118270210208561e+01, // 604
-6.010784439223481e+01, // 605
 3.077858425448244e+02, // 606
 6.929257007056261e+02, // 607
 2.984653305868814e+02, // 608
-6.351276831512137e+02, // 609
-2.689615160495883e+02, // 610
 3.134708140780401e+02, // 611
 4.924433648542910e+02, // 612
-3.094791489648469e+01, // 613
-3.393641704336048e+00, // 614
-1.102157388204757e+02, // 615
 1.436293899423695e+02, // 616
-4.062428270476360e+02, // 617
-1.314457589986538e+02, // 618
 1.194413621647943e+02, // 619
 1.004169408164201e+03, // 620
 1.083398862571992e+02, // 621
-1.595168184290201e+02, // 622
-2.932749395815260e+01, // 623
-1.686279748336820e+01, // 624
-1.894946828374674e+02, // 625
-3.028025448311489e+02, // 626
 4.645457987719102e+02, // 627
-9.582718179191594e+02, // 628
 4.586800910772961e+02, // 629
-8.579900414084199e+01, // 630
 3.642801543052582e+02, // 631
 3.460837927438826e+00, // 632
 2.326131157216161e+02, // 633
 2.335614878256055e+02, // 634
 1.346780228224405e+02, // 635
 1.254112193078151e+02, // 636
 2.856156250715003e-01, // 637
 1.139550540886461e+02, // 638
 1.141610812350877e+02, // 639
-3.659504023940175e-01, // 640
-8.070147392613615e-01, // 641
-1.290416141592268e+02, // 642
-2.086578039734223e+02, // 643
-8.121444349740251e+00, // 644
 1.337463403962308e+02, // 645
-9.690335153925800e+01, // 646
-4.319684237173463e+01, // 647
 2.050681102597557e+01, // 648
-4.506339293519066e+02, // 649
 6.228320359088552e+01, // 650
 4.717281490296572e+01, // 651
 3.351158122952807e+01, // 652
-4.265055339872847e+01, // 653
-1.369880419631458e+02, // 654
-8.926771329181570e+01, // 655
-3.228330693081396e+01, // 656
 3.125532878138061e+01, // 657
-1.615981883773933e+02, // 658
 2.813477402639182e+02, // 659
 3.822462742084146e+01, // 660
 9.991639448215558e+01, // 661
 6.783839880442986e+01, // 662
 2.048348528250254e+02, // 663
-8.348437912997130e+01, // 664
 2.030678822781450e+01, // 665
 8.258001911222037e+01, // 666
 1.466007634277043e+02, // 667
 7.893010581543944e+02, // 668
-1.194400503790063e+02, // 669
 6.681858445360818e+01, // 670
-4.726773896260219e+01, // 671
 5.013962102529787e+02, // 672
 8.607601674333067e+01, // 673
 6.016119673306176e+02, // 674
-7.148928465092846e+00, // 675
 6.064152711213902e+01, // 676
 2.471173407579416e+01, // 677
 4.098013334811909e-01, // 678
-3.616665503501347e+01, // 679
-2.489532874906375e+01, // 680
-8.891675294200966e-01, // 681
-3.799413099293000e+01, // 682
-6.926152054127655e+01, // 683
 1.352444086519573e+02, // 684
-8.205909028598896e+01, // 685
-7.757636631684320e+00, // 686
-1.801324357658820e+02, // 687
-2.072790999931452e+02, // 688
 2.595711841708940e+02, // 689
-2.626996394522333e+01, // 690
 7.043640857535883e+01, // 691
 1.054084527153309e+02, // 692
 4.363813403872821e+01, // 693
 1.328103049954748e+02, // 694
-4.360691269583710e+02, // 695
-4.842947417857398e+01, // 696
-3.710766375224567e+01, // 697
-5.618628230369639e+01, // 698
 4.028625722018445e+01, // 699
-1.153451809540943e+01, // 700
 2.899896081139885e+02, // 701
-2.648055523539025e+01, // 702
-1.635756135876374e+02, // 703
 3.526002011293356e+02, // 704
 6.260438701017105e+01, // 705
-1.178256151994970e+02, // 706
-2.477090228221084e+02, // 707
 2.955263699540606e+02, // 708
-4.794194654223494e+02, // 709
-4.122819692642823e+01, // 710
-7.422016202737505e+01, // 711
 3.845280087151534e+02, // 712
 1.434563997352558e+02, // 713
-1.273786895355677e+03, // 714
-8.197672428140818e+01, // 715
 1.044889675626683e+01, // 716
-2.594753552903632e+02, // 717
 5.682455758540953e+02, // 718
 2.090178678632215e+02, // 719
 6.153623074382520e+01, // 720
 1.157962568844677e+02, // 721
 7.716318542160882e+01, // 722
-1.618072493126122e+02, // 723
-1.709893790554868e+02, // 724
-7.599336835783887e+02, // 725
 1.132832085360454e+02, // 726
-1.984608468318925e+02, // 727
-2.671249764189679e+02, // 728
-1.050522113709704e+03, // 729
 9.669002616869632e+00, // 730
-1.684455006779536e+02, // 731
-2.035479018202778e+02, // 732
 6.199723986620931e+00, // 733
-3.154431782675284e+02, // 734
 1.058576004529692e+02, // 735
 5.847283864300797e+02, // 736
-3.549725704991445e+01, // 737
 1.335238399579943e+01, // 738
 5.896319718629993e+02, // 739
 8.186674918672099e+01, // 740
-7.824859714881145e+00, // 741
-2.011669556812757e+02, // 742
 1.729835225813751e+00, // 743
 1.159543908438835e+02, // 744
-1.502740262256524e+02, // 745
 7.572970725961159e+01, // 746
-2.730827582697162e+02, // 747
-7.782757154052653e+01, // 748
 2.146681025053870e+01, // 749
 2.848353809803719e+02, // 750
 5.558253963238809e+01, // 751
 1.992332732091363e+01, // 752
-2.717606352972363e+01, // 753
 1.948131280099925e+01, // 754
 2.083100021740354e+01, // 755
-1.008463192566674e+02, // 756
 3.069520441084136e+01, // 757
-1.048033764728557e+02, // 758
-8.085716308214799e+01, // 759
-5.800272356397242e+01, // 760
 2.159634893674719e+02, // 761
 2.664985892127254e+01, // 762
 1.351727047458780e+02, // 763
-1.465890728370753e+02, // 764
 5.175224193843444e+01, // 765
 4.394841691763138e+01, // 766
 1.915549592792675e+02, // 767
-3.027295318309572e+02, // 768
-1.230847575072511e+02, // 769
-5.536098709996833e+01, // 770
-5.865290437541286e+00, // 771
 2.002502759440874e+02, // 772
-9.961557632208078e+01, // 773
 9.113025716040437e+01, // 774
 3.630504131772140e+00, // 775
-4.648977371453550e+01, // 776
 2.416671686764419e+02, // 777
-5.025781399395300e+02, // 778
 7.849519765195546e+01, // 779
-9.240656340134491e-01, // 780
-1.394710316930091e+02, // 781
-1.007393112465326e+02, // 782
-8.837332172463588e+00, // 783
 5.395637517827006e+02, // 784
 5.415852013743712e+01, // 785
 8.269210560829288e+00, // 786
-8.625287258710383e+00, // 787
 2.069223863838585e+02, // 788
 2.299209579632790e+02, // 789
-1.333456456555654e+02, // 790
 9.384834115700046e+01, // 791
-4.444763364238143e+02, // 792
 1.364337961310658e+02, // 793
 2.503011475079038e+02, // 794
 1.519738945313279e+02, // 795
-5.792937700749872e+00, // 796
-2.697370519886674e+02, // 797
 4.163121890840901e+02, // 798
-3.743041993021100e+02, // 799
-5.121576346128856e+00, // 800
 4.660312779852590e+01, // 801
-9.448861970373640e+00, // 802
-3.292979094941064e+01, // 803
-4.924833282147465e+01, // 804
-9.098464902779732e+01, // 805
-2.255148870469795e+02, // 806
-1.956593036771320e+02, // 807
-2.641547793622757e+02, // 808
 1.961695493360494e+02, // 809
 1.993624599910206e+00, // 810
-3.393730540548664e+02, // 811
 1.423429473925135e+02, // 812
-3.860182062773337e+00, // 813
-1.829542812824222e+02, // 814
-1.041693760727627e+02, // 815
 4.242726501184443e+02, // 816
 2.851222561351414e+02, // 817
-3.837122668127720e+02, // 818
-8.060771432487027e+01, // 819
 4.623497198893979e+01, // 820
 4.590040776731819e-01, // 821
 5.976562030719321e+01, // 822
 2.579179809483724e+01, // 823
 2.643096933412909e-02, // 824
 2.543666265796348e+01, // 825
-1.887658423594246e-02, // 826
-1.137616458728547e+02, // 827
-2.485033342930738e+02, // 828
-1.069428475437283e+00, // 829
 2.933282592333192e+01, // 830
 4.956245293714383e+01, // 831
 9.772634520060431e+01, // 832
-1.576869697299048e+02, // 833
-8.526410184254370e+01, // 834
-1.019166127957405e+02, // 835
 1.030233967337827e+01, // 836
 4.152488703705850e+01, // 837
 2.032801443369828e+01, // 838
-1.126760528133935e+02, // 839
 3.579273554063957e+01, // 840
 1.263366965045343e+01, // 841
-7.517569463422475e+01, // 842
 6.188119276853463e+02, // 843
 8.365906475805268e+00, // 844
-2.517827192751460e+01, // 845
 3.896280482763352e+00, // 846
 1.681800708034905e+02, // 847
 1.122044616226688e+02, // 848
 2.153073939174307e+01, // 849
 1.543481827556935e-02, // 850
 1.392718666968072e+01, // 851
-7.279889386034182e-02, // 852
 2.323979737932463e+01, // 853
 1.053661507100168e+01, // 854
 1.616419958584345e+02, // 855
-1.385376175638386e+02, // 856
-1.054686292638993e+02, // 857
-2.021600532719876e+02, // 858
-2.934408625673488e+02, // 859
-2.763650861158388e+01, // 860
 2.267440849036536e+01, // 861
-2.027229547776468e+02, // 862
-9.963872374695120e+01, // 863
 3.274829062592844e+02, // 864
-2.603605784787896e+02, // 865
-3.270237244440619e+01, // 866
-1.359609736275077e+02, // 867
-1.106088501125460e+02, // 868
 4.645457886528696e+02, // 869
 1.056268523331892e+03, // 870
 1.512688844218808e+02, // 871
 4.909037413710091e+01, // 872
 1.323175637438483e+02, // 873
 3.201741897466607e+02, // 874
 1.349331008129433e+01, // 875
-1.028346294012907e+02, // 876
 1.609222195773340e+02, // 877
 7.657596569519710e+01, // 878
-4.017490685382514e+01, // 879
-4.775542539195886e+02, // 880
-6.610964038687023e+01, // 881
 2.119653840203537e+03, // 882
 1.953183852998352e+03, // 883
 8.043037221545967e+01, // 884
 2.728162070038053e+02, // 885
 7.297415451268401e+01, // 886
-2.662210448166700e+02, // 887
 6.857911816283409e+01, // 888
 2.480505614377401e+02, // 889
-1.536900825802746e+02, // 890
-2.923720662207502e+02, // 891
-2.641199681814356e-01, // 892
-9.680647362661762e+01, // 893
 2.546053519152277e+02, // 894
 8.839861760369693e+01, // 895
 9.065393488716541e+01, // 896
 1.989247415374844e+00, // 897
 2.262840928884022e+01, // 898
-1.350127265868050e+01, // 899
 1.080613943629697e+02, // 900
 9.150831778951326e+01, // 901
 3.514127935145757e+01, // 902
 1.141567415424944e+02, // 903
 3.091934591187341e+02, // 904
-6.253530583409945e+01, // 905
 5.658310819709055e+00, // 906
-2.152163930316658e+02, // 907
-2.205119423084873e+01, // 908
-5.611678424123192e+01, // 909
-8.297007324529620e+00, // 910
-5.723785915152487e+00, // 911
 1.701766512076007e+02, // 912
 2.576083349853322e+02, // 913
-3.791439173522279e+01, // 914
-1.616200763375622e+02, // 915
 8.181117369039158e+01, // 916
-1.634947638336631e+02, // 917
-1.023450388036669e+02, // 918
 4.086382510442789e+01, // 919
-2.186335174230369e+02, // 920
-1.120049416300434e+02, // 921
-3.547178277664236e+01, // 922
-2.033358478301910e+02, // 923
 7.046285222115536e+01, // 924
 3.229620385756101e+02, // 925
 1.291974442276382e+02, // 926
 6.231008162432747e+02, // 927
 3.326421152954794e+02, // 928
 2.021316285876889e+02, // 929
 1.709063444482635e+02, // 930
 1.048186698233212e+02, // 931
 1.469689979240223e+02, // 932
-6.720265152771610e+01, // 933
 3.642901870626988e+00, // 934
-2.908197223636149e+02, // 935
 2.519325625916446e+02, // 936
 5.080408906746530e+00, // 937
-9.737000910668266e+01, // 938
-7.878994057188126e+01, // 939
 8.538284560441760e+01, // 940
-1.355936242669253e+01, // 941
 8.098072120800263e+02, // 942
 1.154030489811840e+03, // 943
-2.452932339518815e+02, // 944
 8.965292156895381e+01, // 945
-1.944537346072658e+01, // 946
 3.440893026049677e+02, // 947
 5.724288154240768e+02, // 948
 8.493175873621259e+01, // 949
 4.784888470182066e+01, // 950
 5.129035576756011e+01, // 951
 2.257866644150775e+00, // 952
 1.218926777076382e+00, // 953
-3.366044836090475e-03, // 954
 2.500772101705775e+02, // 955
 1.490471702781856e+02, // 956
 3.813681869357914e+01, // 957
 5.587503886147421e-01, // 958
 6.559089773914150e+00, // 959
-7.280295532960592e+01, // 960
 2.999363878062402e+00, // 961
 1.905290805077184e+00, // 962
 2.689738181696958e-03, // 963
 1.475698807527274e+00, // 964
-5.400120548054011e-03, // 965
-5.856036381543734e+01, // 966
-7.466333318161814e+01, // 967
-1.410484600880401e+02, // 968
 1.890809963291293e-01, // 969
 9.322524177136573e+00, // 970
-1.058227379834338e+02, // 971
 8.095391617749773e-01, // 972
-3.593616800769065e+01, // 973
-9.456712229617580e+01, // 974
-1.271879392917515e+02, // 975
-1.056770637869856e+02, // 976
 3.854288213948202e-01, // 977
-3.767873796691350e+01, // 978
 5.298387851148630e-01, // 979
-8.037854356391128e+01, // 980
-3.700079168055471e+01, // 981
-3.313877841830263e+01, // 982
-9.791466768782570e+01, // 983
-1.416981602098307e+02, // 984
 9.297968056829697e-01, // 985
-3.357420710326281e+01, // 986
-2.114797107826883e+02, // 987
-2.390826030589256e-01, // 988
-6.781870407397066e+01, // 989
-1.465452513174128e+02, // 990
-1.037099072844005e+02, // 991
 1.607141611586006e+02, // 992
 1.134763764459052e+00, // 993
 9.993420662085170e+01, // 994
 9.812833672381898e+01, // 995
 6.218954429675562e+01, // 996
-6.791288563899583e+01, // 997
 5.103122673051875e-01, // 998
-1.429860422198564e+02, // 999
 2.083076430850956e-02, // 1000
-8.091727870559332e+01, // 1001
-4.743371563216166e+01, // 1002
 2.289711325145655e+02, // 1003
 8.363527685222461e+01, // 1004
 2.494417047915242e+02, // 1005
 9.366643271284944e+01, // 1006
-1.515052830328407e+01, // 1007
-1.430943247934581e+01, // 1008
-4.664358712619908e+01, // 1009
 2.001263899016383e+00, // 1010
 1.168776346005158e+02, // 1011
 9.106507376112974e+00, // 1012
 2.154729444987463e+00, // 1013
-9.849583623545779e+01, // 1014
-1.278884103832939e+02, // 1015
-1.598649827435965e+02, // 1016
 6.534104407774008e+01, // 1017
-1.949630114244436e+02, // 1018
 1.096527429838266e+02, // 1019
 1.406833286454741e+01, // 1020
-9.552609284911424e+01, // 1021
 2.960078798125223e-01, // 1022
-7.815389654327637e+01, // 1023
 2.451200389530512e-01, // 1024
-7.280362639927027e+01, // 1025
 1.187711426926927e-01, // 1026
-6.198350824921858e+01, // 1027
-2.257199471376295e+01, // 1028
-7.004560027896123e+00, // 1029
 4.431199071672469e+01, // 1030
-3.995901271204551e+01, // 1031
 2.025555632060167e+00, // 1032
-8.299795173756121e+01, // 1033
-3.057629331658385e+02, // 1034
-2.362969216195194e+02, // 1035
-8.388550870467013e+01, // 1036
 1.713336668879226e+02, // 1037
 2.093627553122144e+02, // 1038
 1.384231013042848e+02, // 1039
 1.578119487651454e-01, // 1040
 1.328572951902611e+02, // 1041
-1.192367839811673e-01, // 1042
 6.939751193497146e+01, // 1043
-1.049583768838877e+02, // 1044
-2.318633764457365e+02, // 1045
 4.494144353217747e+01, // 1046
-6.330300596145517e+01, // 1047
-3.170540349745034e+02, // 1048
 3.322022358336895e+02, // 1049
 1.513020505216568e+02, // 1050
 3.705474463138562e+01, // 1051
 1.422171676943055e+01, // 1052
 1.645670601447553e+02, // 1053
-1.730580143977255e+01, // 1054
 1.719238618350258e+01, // 1055
 3.149488111224225e+02, // 1056
 7.100833322923371e+01, // 1057
-2.102569282062714e+00, // 1058
-8.776290259241917e+01, // 1059
-3.086597288396325e+02, // 1060
-4.670510829273054e+01, // 1061
-1.433904710972018e+02, // 1062
 1.117875580388317e+02, // 1063
-3.115018780364193e+01, // 1064
 2.556351473821618e+01, // 1065
-4.854397986046041e+02, // 1066
 6.088548331320678e+01, // 1067
-1.682658036375701e+02, // 1068
-2.636750304687854e+02, // 1069
 2.333465283299905e+02, // 1070
 2.040408802461952e+02, // 1071
 3.708082275078710e+01, // 1072
 1.018795846325803e+02, // 1073
 1.928552251164243e+01, // 1074
 3.239858735125246e+01, // 1075
 2.676085269129110e+02, // 1076
 1.786778371702901e+02, // 1077
 4.959254127782724e+01, // 1078
-5.076782596064187e+01, // 1079
 1.620025265964809e+02, // 1080
-3.012945484267810e+01, // 1081
-3.055587991250038e+01, // 1082
 1.786653478360953e+02, // 1083
-6.745426864463627e+01, // 1084
-4.917190718480749e+01, // 1085
-6.081172056066193e+01, // 1086
-2.229221332250890e+02, // 1087
 2.249862623586424e+01, // 1088
-4.355796204054511e+01, // 1089
-6.918209134899784e+01, // 1090
-3.557551658866272e+02, // 1091
-1.923864403879129e+01, // 1092
-1.441377772021342e+02, // 1093
-1.436290248864072e+02, // 1094
-2.192371796436579e+01, // 1095
 1.082351954653423e+02, // 1096
 1.989715771486069e+02, // 1097
-1.575810959383425e+02, // 1098
-1.805969421829489e+02, // 1099
 8.984723324614466e+02, // 1100
 5.806703342296659e+02, // 1101
 6.359149250082321e-01, // 1102
 5.666288308237368e+02, // 1103
-4.050916881149930e-01, // 1104
-1.847180333897176e+02, // 1105
 8.110877831821463e+01, // 1106
 1.959748388225103e+02, // 1107
 1.912932554699908e+02, // 1108
-2.315519087199365e+01, // 1109
-3.246569024173722e+02, // 1110
 2.120850027145839e+02, // 1111
-7.195367905732680e+01, // 1112
 1.526568489029964e+02, // 1113
-6.045913268860706e+01, // 1114
 6.079398284779486e+02, // 1115
-9.089616633608782e+01, // 1116
 6.600647840561389e+01, // 1117
-7.568117228962680e+01, // 1118
 2.036326996876174e+02, // 1119
-9.829482433049751e+01, // 1120
-6.593177579258177e+01, // 1121
 1.387854348793928e+02, // 1122
 7.872258700023771e+01, // 1123
-3.550461150056411e+02, // 1124
 1.591905203149350e+02, // 1125
-5.393697085470592e+01, // 1126
-2.575260868311113e+01, // 1127
-9.892581703875975e+01, // 1128
 1.750834157408007e+02, // 1129
-3.170608369713416e+02, // 1130
 3.320675321093140e+01, // 1131
 3.543040543791129e+02, // 1132
 1.527190907971383e+02, // 1133
 2.475669126611468e+02, // 1134
-4.301381480943443e+00, // 1135
 2.659239282758317e+01, // 1136
 4.672164961560176e+01, // 1137
-1.597188639785293e+02, // 1138
 1.007642214217297e+02, // 1139
-1.319385289895205e+01, // 1140
-2.516923355867251e+01, // 1141
 2.764356009498134e+02, // 1142
-2.531548633350027e+01, // 1143
 9.564204000574216e+01, // 1144
 1.763430344678988e+02, // 1145
 9.471782087263398e-01, // 1146
 1.757015149773515e+02, // 1147
 6.253363098815754e+01, // 1148
 1.221474060573705e+02, // 1149
 8.764116232123472e+01, // 1150
-1.513395903424437e+02, // 1151
 4.807131512095127e+01, // 1152
-9.038553968648125e+01, // 1153
-3.309322814484569e+02, // 1154
-2.591182671330873e+02, // 1155
-3.541783057615153e+02, // 1156
-1.703105057505226e+01, // 1157
 9.189558847916450e+01, // 1158
 6.729717887552819e+01, // 1159
 7.641628746388376e+02, // 1160
 1.616193366010608e+02, // 1161
-2.107313843962473e+02, // 1162
 4.313342342380265e+02, // 1163
-7.364578462755708e+01, // 1164
 7.261753951094445e+01, // 1165
 1.292762833138370e+02, // 1166
-2.376359484524767e+01, // 1167
 1.710125401003312e+02, // 1168
-1.773952515308396e+02, // 1169
 2.788379078600353e+01, // 1170
 7.825281732771914e+01, // 1171
-1.128222805595669e+02, // 1172
-1.135239226536850e+02, // 1173
 9.506307322506144e+01, // 1174
-9.451366681119568e+01, // 1175
 1.358534609905517e+00, // 1176
-1.096310441054451e+02, // 1177
-1.390634182321940e+02, // 1178
-3.292329564779187e+02, // 1179
-3.023547839550776e+02, // 1180
-1.438788951042639e+02, // 1181
-5.621803649222635e+02; // 1182

}

netcdf mbnrg_1b_A1B3C1D2_fit {
  // global attributes 
  :name = " mbnrg_1b_A1B3C1D2_fit";
  :k_x_intra_A_B_1 =  1.002770900240316e+00; // A^(-1))
  :k_x_intra_A_C_1 =  1.474647851755247e+00; // A^(-1))
  :k_x_intra_A_D_1 =  2.579994050104364e-01; // A^(-1))
  :k_x_intra_B_B_1 =  4.972427481128774e-01; // A^(-1))
  :k_x_intra_B_C_1 =  4.058760621697250e-01; // A^(-1))
  :k_x_intra_B_D_1 =  4.768645823601143e-01; // A^(-1))
  :k_x_intra_C_D_1 =  1.213760623498014e+00; // A^(-1))
  :k_x_intra_D_D_1 =  6.313929230907642e-01; // A^(-1))
  :ri =  0.000000000000000e+00; // A
  :ro =  0.000000000000000e+00; // A
  dimensions:
  poly = 353;
  variables:
    double poly(poly);
data:
poly =
 7.890961170423259e+01, // 0
 7.692882665149973e+02, // 1
-3.600194922660839e+03, // 2
 8.267477678959024e+02, // 3
-1.807854642917589e+03, // 4
 4.322829515378949e+03, // 5
-3.913834078247157e+02, // 6
-6.184969416913523e+02, // 7
-9.241088157177689e+02, // 8
 6.170532577244861e+02, // 9
 1.509920721342151e+02, // 10
 4.465317489748783e+03, // 11
 8.244626921659627e+02, // 12
 2.745059023001278e+02, // 13
 3.738645157237743e+02, // 14
-2.268522941966353e+02, // 15
-3.642863662661039e+02, // 16
 2.974481701063529e+02, // 17
-1.058858234081164e+03, // 18
-8.817222443276601e+02, // 19
 4.223364729741796e+02, // 20
 8.263965616111980e+02, // 21
 2.062577714230351e+00, // 22
 3.966148287104229e+02, // 23
 1.193453834640986e+02, // 24
-2.633412401065461e+02, // 25
 1.706432419274805e+02, // 26
-7.716214752335839e+02, // 27
-7.990635770570734e+01, // 28
-3.574872200238735e+01, // 29
 2.281684357508506e+03, // 30
 1.180022140684204e+03, // 31
 1.320598253814275e+02, // 32
 9.985765232005817e+02, // 33
-1.071925675887201e+03, // 34
-7.163712918345410e+02, // 35
-1.886295238161705e+02, // 36
-2.814451284672895e+02, // 37
 1.398531882254090e+02, // 38
-2.504214572729120e+02, // 39
 1.093663258465553e+02, // 40
-1.138066065145470e+03, // 41
 2.649565100723573e+03, // 42
 1.024308026243941e+03, // 43
-2.242087051243618e+02, // 44
-3.857098284019844e+01, // 45
 1.417376790734048e+02, // 46
-1.682472756533483e+01, // 47
-5.134503181331361e+02, // 48
-2.196087714094973e+02, // 49
 2.712139958210859e+02, // 50
 5.558313093385980e+02, // 51
 5.196774611182133e+02, // 52
-8.999804562495742e+02, // 53
 2.623251242948912e+03, // 54
-2.517115702270120e+03, // 55
-1.553674861126279e+03, // 56
 7.159735954195894e+02, // 57
-9.228170016674746e+02, // 58
-6.017214029277322e+02, // 59
 8.926164862829594e+02, // 60
-3.569063144032315e+03, // 61
-1.286932585937038e+03, // 62
-8.211204182799294e+02, // 63
 3.722325585987615e+00, // 64
 5.291353269994223e+02, // 65
-1.013950307670441e+03, // 66
-4.380477420318887e+02, // 67
 1.259194002670791e+03, // 68
 1.397578088340010e+03, // 69
 2.893228842373919e+03, // 70
-2.255540263585223e+03, // 71
-8.344922073772988e+02, // 72
-1.931285374493160e+02, // 73
 6.127697245208377e+02, // 74
-2.890540811426001e+02, // 75
 1.866632415187280e+03, // 76
-1.302635477068233e+03, // 77
-1.603925848182814e+03, // 78
 1.479024865344926e+03, // 79
 1.609530791481580e+02, // 80
 2.635517616778226e+02, // 81
 8.612222610230393e+01, // 82
-2.250186370844195e+02, // 83
 5.584576239407840e+00, // 84
 1.707880084295927e+02, // 85
-3.143184890689525e+01, // 86
-1.405964901873654e+01, // 87
-5.349922421466832e+02, // 88
 4.144502210242542e+02, // 89
 2.698246203908801e+02, // 90
 1.818387488272886e+02, // 91
 1.435947463965109e+02, // 92
-6.626285894197811e+02, // 93
 1.514589323192409e+02, // 94
-7.057836221843399e+02, // 95
-1.481579361140836e+03, // 96
-3.865736917398165e+02, // 97
 8.514324505534168e+01, // 98
 1.726174688861166e+02, // 99
-3.302837984670356e+02, // 100
 3.551803716045775e+02, // 101
-1.094086273193941e+03, // 102
 1.125473925974490e+03, // 103
-4.960730708009792e+01, // 104
 2.548785087310909e+03, // 105
-1.221827461918868e+03, // 106
 8.939630409843642e+02, // 107
 3.549556249112364e+02, // 108
-7.790864486703174e+01, // 109
-1.901431971459646e+02, // 110
 9.766685856982740e+02, // 111
 5.925904992874161e+01, // 112
-2.564907919443181e+03, // 113
-2.845505029061504e+03, // 114
 4.883662993878351e+02, // 115
 2.716028032006936e+03, // 116
-8.507623961397924e+02, // 117
-1.353305119027594e+02, // 118
-9.257628524798442e+02, // 119
 1.120683645974798e+03, // 120
 1.922457189413646e+03, // 121
-1.868374049144599e+03, // 122
-2.165320487012457e+03, // 123
-5.555729865074378e+03, // 124
-1.003952566793386e+03, // 125
-2.560890696045740e+02, // 126
 4.201256302012998e+02, // 127
-7.640858738006515e+02, // 128
-1.596208545566165e+03, // 129
-1.258602275878287e+02, // 130
 7.561148579101230e+02, // 131
 1.522124168356052e+03, // 132
-4.548986096598542e+02, // 133
-3.704097909306405e+02, // 134
-6.416348028544812e+02, // 135
 9.480199607456601e+02, // 136
 1.874763778215718e+02, // 137
-1.017256160134526e+03, // 138
-2.556272309380266e+01, // 139
-8.534191599212892e+02, // 140
-1.143616828299137e+03, // 141
-7.647156791675917e+00, // 142
 2.521357745690285e+02, // 143
-1.579046269741806e+03, // 144
-2.762472120312184e+03, // 145
-4.934664834790877e+02, // 146
-5.027447292770917e+02, // 147
 6.979791141460545e+02, // 148
 9.841671968842967e+02, // 149
 4.914918816176747e+02, // 150
 1.743936596749943e+03, // 151
-5.806721870358635e+01, // 152
 2.897857564670422e+03, // 153
 3.599540363397664e+02, // 154
-9.390067822181654e+02, // 155
 1.060093785062037e+03, // 156
-3.277030180458126e+03, // 157
-5.599886246753312e+02, // 158
 6.213751013489513e+02, // 159
 2.684739684410868e+02, // 160
-1.843787737462930e+03, // 161
-1.010444431962834e+03, // 162
 1.979834521940816e+03, // 163
-1.450568515514235e+03, // 164
 1.555811848037474e+03, // 165
 4.165668278344671e+01, // 166
 5.827057493358168e+02, // 167
-2.109006602167225e+02, // 168
 1.952867779287844e+02, // 169
 1.038706731448365e+03, // 170
-1.060214063197115e+03, // 171
 5.815805231032742e+01, // 172
-7.812048866945174e+02, // 173
-5.119909983701285e+02, // 174
 3.271615556866931e+01, // 175
 3.631474955804622e+02, // 176
-7.823773266021198e+02, // 177
 2.317155133874491e+02, // 178
 2.052289602963436e+02, // 179
-1.138552931737795e+03, // 180
-1.420482965975623e+03, // 181
-6.796405248328300e+02, // 182
 1.352543899805003e+03, // 183
-8.710264669516251e+02, // 184
 2.424475202437056e+02, // 185
 1.933798984420329e+02, // 186
 9.515242778382693e+02, // 187
 4.434122500399367e+02, // 188
 1.965171607525363e+03, // 189
 3.635511776293489e+02, // 190
-1.975205251404725e+03, // 191
 1.897950654841097e+03, // 192
 2.161367479321688e+02, // 193
 2.444047204787014e+02, // 194
 2.196122244510083e+02, // 195
-1.430202313789307e+01, // 196
 2.218675673809987e+02, // 197
 1.445537631819407e+01, // 198
-1.918192274397658e+02, // 199
 2.694278568711800e+02, // 200
-8.587203781792186e+01, // 201
-1.557337487475026e+02, // 202
-8.728719620536367e+02, // 203
-2.026917493734558e+02, // 204
 3.507856462757139e+02, // 205
-5.478061335090471e+02, // 206
-1.138839342361392e+03, // 207
 1.515769412266209e+03, // 208
 1.334040366667227e+01, // 209
 1.315812670772784e+03, // 210
 4.689662903821439e+02, // 211
 5.634047719093767e+02, // 212
 1.105414894379277e+03, // 213
-4.787527694836887e+02, // 214
 5.144126863613496e+02, // 215
 1.136084025444600e+03, // 216
 2.130110460527740e+03, // 217
 5.365238995522213e+02, // 218
 2.736893229860449e+02, // 219
-1.932251847654015e+02, // 220
 5.548795014130020e+02, // 221
 2.276431531992947e+02, // 222
-3.774913712810549e+02, // 223
 1.566341351338087e+01, // 224
 7.119791580705275e+02, // 225
 4.379440419127278e+02, // 226
-1.098379775235203e+03, // 227
-2.219801012099581e+01, // 228
-2.649248453203400e+02, // 229
-5.817943863705868e+02, // 230
-1.630460997900339e+03, // 231
 1.894436158257042e+03, // 232
-3.449330470654352e+02, // 233
-2.258323033525279e+02, // 234
-5.342133461103419e+02, // 235
 4.992231598234389e+02, // 236
 4.125829478348076e+02, // 237
 2.281730850601871e+02, // 238
 4.060943124975988e+02, // 239
 1.255585196480816e+03, // 240
 1.284827439516299e+03, // 241
 5.803982738566305e+02, // 242
 8.023812037086495e+02, // 243
 5.414684567953237e+02, // 244
-1.930152353106872e+02, // 245
 3.369132106487078e+02, // 246
 5.391378073243434e+02, // 247
-5.430089918501930e+02, // 248
 1.358831009275251e+02, // 249
-1.488514024143615e+02, // 250
 1.945979755178894e+01, // 251
-3.308117694301047e+01, // 252
-4.346469475374261e+02, // 253
 2.866203907850135e+02, // 254
-2.732099668071974e+02, // 255
-9.068253257852315e+02, // 256
-2.333678154805375e+01, // 257
 8.709098412793174e+02, // 258
-6.795505735066124e+02, // 259
 2.002113946633959e+02, // 260
 7.926428480868805e+01, // 261
 5.266944799922943e+01, // 262
 7.896828851499199e+02, // 263
 3.227960461043137e+02, // 264
-4.373126308154611e+02, // 265
-4.930665308208883e+02, // 266
 3.997922219304219e+02, // 267
 2.062549930613451e+02, // 268
 2.934450215879244e+02, // 269
 7.546048595317566e+02, // 270
 4.482618595649964e+02, // 271
-3.112486357072370e+02, // 272
 2.785649697628627e+02, // 273
-4.592726375073193e+02, // 274
-5.754039328177922e+02, // 275
 1.670976695608693e+03, // 276
 6.967566610762668e+01, // 277
-6.522936044872511e+02, // 278
-2.991607760547091e+02, // 279
 7.497679523532253e+01, // 280
 8.065868754337703e+02, // 281
-1.489010245152553e+03, // 282
-8.807375474900261e+02, // 283
-3.302896771015253e+02, // 284
-3.405470712647502e+01, // 285
 1.606760401902206e+02, // 286
-6.663972767574007e+02, // 287
 1.024056476922640e+02, // 288
 1.888349500109766e+03, // 289
 2.743729157907807e+03, // 290
-9.422421391533589e+02, // 291
 5.908035942690807e+01, // 292
 7.837133837825950e+02, // 293
-1.671732522252044e+01, // 294
 1.368146682877980e+03, // 295
-5.361967839405677e+02, // 296
-1.019285071375023e+02, // 297
-1.912810653927410e+03, // 298
 7.060520775926104e+02, // 299
-3.943378497834835e+02, // 300
 8.622444085406940e+01, // 301
 1.382664274417756e+03, // 302
-9.156337846061219e+02, // 303
-2.538928328998821e+02, // 304
 1.050660200103816e+02, // 305
-1.166703449320033e+03, // 306
-4.973478539999977e+01, // 307
 1.236077402496876e+03, // 308
 3.263582954945890e+02, // 309
 3.151162415958993e+02, // 310
-2.553353445031327e+02, // 311
-2.314146265117134e+02, // 312
-1.398060751795938e+03, // 313
 4.304071670968367e+02, // 314
-7.689950628017745e+02, // 315
 1.135739741533998e+03, // 316
-4.515219736840731e+02, // 317
-3.052648713963722e+02, // 318
-6.509505046072293e+02, // 319
-9.138768408643684e+02, // 320
 1.584046003272575e+02, // 321
-1.144412009682541e+02, // 322
-6.595547928684055e+02, // 323
 1.026181210759939e+01, // 324
 8.048601470590920e+02, // 325
-1.680935719281379e+03, // 326
 3.422702966597776e+02, // 327
-3.717380806230411e+02, // 328
 1.677858569832690e+02, // 329
-1.835467111971880e+02, // 330
-5.146657972956500e+02, // 331
-5.160599137812380e+02, // 332
 2.554885292464364e+02, // 333
-2.046519573659203e+02, // 334
 4.344899959447337e+02, // 335
-5.329339472711199e+01, // 336
-2.912005291498753e+01, // 337
-2.634108901920640e+02, // 338
-9.151076753824015e+01, // 339
-1.057613233378803e+03, // 340
 6.656089745954557e+01, // 341
 3.345051875132287e+02, // 342
-8.159766511977637e+01, // 343
 8.056747574709733e+02, // 344
 6.784161539965862e+01, // 345
-2.336435221085117e+02, // 346
 5.114860819120543e+02, // 347
 3.075917412646961e+02, // 348
-5.838808467629118e+02, // 349
 8.167758405856246e+00, // 350
-9.913427282368021e+02, // 351
 4.068710212404188e+03; // 352

}

netcdf mbnrg_2b_A1B3C1D2_E1F2_fit {
  // global attributes 
  :name = " mbnrg_2b_A1B3C1D2_E1F2_fit";
  :k_x_intra_A_B_1 =  1.212673330778570e+00; // A^(-1))
  :k_x_intra_A_C_1 =  2.498319716890491e+00; // A^(-1))
  :k_x_intra_A_D_1 =  2.684397328963688e+00; // A^(-1))
  :k_x_inter_A_E_0 =  2.430938657573861e+00; // A^(-1))
  :k_x_inter_A_F_0 =  3.471279829494320e+00; // A^(-1))
  :k_x_intra_B_B_1 =  2.674503866897199e+00; // A^(-1))
  :k_x_intra_B_C_1 =  3.733797571032214e+00; // A^(-1))
  :k_x_intra_B_D_1 =  1.696746596925308e+00; // A^(-1))
  :k_x_inter_B_E_0 =  2.452595534013862e+00; // A^(-1))
  :k_x_inter_B_F_0 =  3.124693258723567e+00; // A^(-1))
  :k_x_intra_C_D_1 =  2.188576351939037e+00; // A^(-1))
  :k_x_inter_C_E_0 =  1.582100203531841e+00; // A^(-1))
  :k_x_inter_C_F_0 =  1.426599549328256e+00; // A^(-1))
  :k_x_intra_D_D_1 =  1.645825476220728e+00; // A^(-1))
  :k_x_inter_D_E_0 =  3.526096316765107e+00; // A^(-1))
  :k_x_inter_D_F_0 =  3.591635413743386e+00; // A^(-1))
  :k_x_intra_E_F_1 =  2.353729987216056e+00; // A^(-1))
  :k_x_intra_F_F_1 =  1.445692745244919e+00; // A^(-1))
  :ri =  6.000000000000000e+00; // A
  :ro =  7.000000000000000e+00; // A
  dimensions:
  poly = 1183;
  variables:
    double poly(poly);
data:
poly =
 0.000000000000000e+00, // 0
 0.000000000000000e+00, // 1
 0.000000000000000e+00, // 2
 0.000000000000000e+00, // 3
 0.000000000000000e+00, // 4
 0.000000000000000e+00, // 5
 0.000000000000000e+00, // 6
 0.000000000000000e+00, // 7
 0.000000000000000e+00, // 8
 0.000000000000000e+00, // 9
 0.000000000000000e+00, // 10
 0.000000000000000e+00, // 11
 0.000000000000000e+00, // 12
 0.000000000000000e+00, // 13
 0.000000000000000e+00, // 14
 0.000000000000000e+00, // 15
 0.000000000000000e+00, // 16
 0.000000000000000e+00, // 17
 0.000000000000000e+00, // 18
 0.000000000000000e+00, // 19
 0.000000000000000e+00, // 20
 0.000000000000000e+00, // 21
 0.000000000000000e+00, // 22
 0.000000000000000e+00, // 23
 0.000000000000000e+00, // 24
 0.000000000000000e+00, // 25
 0.000000000000000e+00, // 26
 0.000000000000000e+00, // 27
 0.000000000000000e+00, // 28
 0.000000000000000e+00, // 29
 0.000000000000000e+00, // 30
 0.000000000000000e+00, // 31
 0.000000000000000e+00, // 32
 0.000000000000000e+00, // 33
 0.000000000000000e+00, // 34
 0.000000000000000e+00, // 35
 0.000000000000000e+00, // 36
 0.000000000000000e+00, // 37
 0.000000000000000e+00, // 38
 0.000000000000000e+00, // 39
 0.000000000000000e+00, // 40
 0.000000000000000e+00, // 41
 0.000000000000000e+00, // 42
 0.000000000000000e+00, // 43
 0.000000000000000e+00, // 44
 0.000000000000000e+00, // 45
 0.000000000000000e+00, // 46
 0.000000000000000e+00, // 47
 0.000000000000000e+00, // 48
 0.000000000000000e+00, // 49
 0.000000000000000e+00, // 50
 0.000000000000000e+00, // 51
 0.000000000000000e+00, // 52
 0.000000000000000e+00, // 53
 0.000000000000000e+00, // 54
 0.000000000000000e+00, // 55
 0.000000000000000e+00, // 56
 0.000000000000000e+00, // 57
 0.000000000000000e+00, // 58
 0.000000000000000e+00, // 59
 0.000000000000000e+00, // 60
 0.000000000000000e+00, // 61
 0.000000000000000e+00, // 62
 0.000000000000000e+00, // 63
 0.000000000000000e+00, // 64
 0.000000000000000e+00, // 65
 0.000000000000000e+00, // 66
 0.000000000000000e+00, // 67
 0.000000000000000e+00, // 68
 0.000000000000000e+00, // 69
 0.000000000000000e+00, // 70
 0.000000000000000e+00, // 71
 0.000000000000000e+00, // 72
 0.000000000000000e+00, // 73
 0.000000000000000e+00, // 74
 0.000000000000000e+00, // 75
 0.000000000000000e+00, // 76
 0.000000000000000e+00, // 77
 0.000000000000000e+00, // 78
 0.000000000000000e+00, // 79
 0.000000000000000e+00, // 80
 0.000000000000000e+00, // 81
 0.000000000000000e+00, // 82
 0.000000000000000e+00, // 83
 0.000000000000000e+00, // 84
 0.000000000000000e+00, // 85
 0.000000000000000e+00, // 86
 0.000000000000000e+00, // 87
 0.000000000000000e+00, // 88
 0.000000000000000e+00, // 89
 0.000000000000000e+00, // 90
 0.000000000000000e+00, // 91
 0.000000000000000e+00, // 92
 0.000000000000000e+00, // 93
 0.000000000000000e+00, // 94
 0.000000000000000e+00, // 95
 0.000000000000000e+00, // 96
 0.000000000000000e+00, // 97
 0.000000000000000e+00, // 98
 0.000000000000000e+00, // 99
 0.000000000000000e+00, // 100
 0.000000000000000e+00, // 101
 0.000000000000000e+00, // 102
 0.000000000000000e+00, // 103
 0.000000000000000e+00, // 104
 0.000000000000000e+00, // 105
 0.000000000000000e+00, // 106
 0.000000000000000e+00, // 107
 0.000000000000000e+00, // 108
 0.000000000000000e+00, // 109
 0.000000000000000e+00, // 110
 0.000000000000000e+00, // 111
 0.000000000000000e+00, // 112
 0.000000000000000e+00, // 113
 0.000000000000000e+00, // 114
 0.000000000000000e+00, // 115
 0.000000000000000e+00, // 116
 0.000000000000000e+00, // 117
 0.000000000000000e+00, // 118
 0.000000000000000e+00, // 119
 0.000000000000000e+00, // 120
 0.000000000000000e+00, // 121
 0.000000000000000e+00, // 122
 0.000000000000000e+00, // 123
 0.000000000000000e+00, // 124
 0.000000000000000e+00, // 125
 0.000000000000000e+00, // 126
 0.000000000000000e+00, // 127
 0.000000000000000e+00, // 128
 0.000000000000000e+00, // 129
 0.000000000000000e+00, // 130
 0.000000000000000e+00, // 131
 0.000000000000000e+00, // 132
 0.000000000000000e+00, // 133
 0.000000000000000e+00, // 134
 0.000000000000000e+00, // 135
 0.000000000000000e+00, // 136
 0.000000000000000e+00, // 137
 0.000000000000000e+00, // 138
 0.000000000000000e+00, // 139
 0.000000000000000e+00, // 140
 0.000000000000000e+00, // 141
 0.000000000000000e+00, // 142
 0.000000000000000e+00, // 143
 0.000000000000000e+00, // 144
 0.000000000000000e+00, // 145
 0.000000000000000e+00, // 146
 0.000000000000000e+00, // 147
 0.000000000000000e+00, // 148
 0.000000000000000e+00, // 149
 0.000000000000000e+00, // 150
 0.000000000000000e+00, // 151
 0.000000000000000e+00, // 152
 0.000000000000000e+00, // 153
 0.000000000000000e+00, // 154
 0.000000000000000e+00, // 155
 0.000000000000000e+00, // 156
 0.000000000000000e+00, // 157
 0.000000000000000e+00, // 158
 0.000000000000000e+00, // 159
 0.000000000000000e+00, // 160
 0.000000000000000e+00, // 161
 0.000000000000000e+00, // 162
 0.000000000000000e+00, // 163
 0.000000000000000e+00, // 164
 0.000000000000000e+00, // 165
 0.000000000000000e+00, // 166
 0.000000000000000e+00, // 167
 0.000000000000000e+00, // 168
 0.000000000000000e+00, // 169
 0.000000000000000e+00, // 170
 0.000000000000000e+00, // 171
 0.000000000000000e+00, // 172
 0.000000000000000e+00, // 173
 0.000000000000000e+00, // 174
 0.000000000000000e+00, // 175
 0.000000000000000e+00, // 176
 0.000000000000000e+00, // 177
 0.000000000000000e+00, // 178
 0.000000000000000e+00, // 179
 0.000000000000000e+00, // 180
 0.000000000000000e+00, // 181
 0.000000000000000e+00, // 182
 0.000000000000000e+00, // 183
 0.000000000000000e+00, // 184
 0.000000000000000e+00, // 185
 0.000000000000000e+00, // 186
 0.000000000000000e+00, // 187
 0.000000000000000e+00, // 188
 0.000000000000000e+00, // 189
 0.000000000000000e+00, // 190
 0.000000000000000e+00, // 191
 0.000000000000000e+00, // 192
 0.000000000000000e+00, // 193
 0.000000000000000e+00, // 194
 0.000000000000000e+00, // 195
 0.000000000000000e+00, // 196
 0.000000000000000e+00, // 197
 0.000000000000000e+00, // 198
 0.000000000000000e+00, // 199
 0.000000000000000e+00, // 200
 0.000000000000000e+00, // 201
 0.000000000000000e+00, // 202
 0.000000000000000e+00, // 203
 0.000000000000000e+00, // 204
 0.000000000000000e+00, // 205
 0.000000000000000e+00, // 206
 0.000000000000000e+00, // 207
 0.000000000000000e+00, // 208
 0.000000000000000e+00, // 209
 0.000000000000000e+00, // 210
 0.000000000000000e+00, // 211
 0.000000000000000e+00, // 212
 0.000000000000000e+00, // 213
 0.000000000000000e+00, // 214
 0.000000000000000e+00, // 215
 0.000000000000000e+00, // 216
 0.000000000000000e+00, // 217
 0.000000000000000e+00, // 218
 0.000000000000000e+00, // 219
 0.000000000000000e+00, // 220
 0.000000000000000e+00, // 221
 0.000000000000000e+00, // 222
 0.000000000000000e+00, // 223
 0.000000000000000e+00, // 224
 0.000000000000000e+00, // 225
 0.000000000000000e+00, // 226
 0.000000000000000e+00, // 227
 0.000000000000000e+00, // 228
 0.000000000000000e+00, // 229
 0.000000000000000e+00, // 230
 0.000000000000000e+00, // 231
 0.000000000000000e+00, // 232
 0.000000000000000e+00, // 233
 0.000000000000000e+00, // 234
 0.000000000000000e+00, // 235
 0.000000000000000e+00, // 236
 0.000000000000000e+00, // 237
 0.000000000000000e+00, // 238
 0.000000000000000e+00, // 239
 0.000000000000000e+00, // 240
 0.000000000000000e+00, // 241
 0.000000000000000e+00, // 242
 0.000000000000000e+00, // 243
 0.000000000000000e+00, // 244
 0.000000000000000e+00, // 245
 0.000000000000000e+00, // 246
 0.000000000000000e+00, // 247
 0.000000000000000e+00, // 248
 0.000000000000000e+00, // 249
 0.000000000000000e+00, // 250
 0.000000000000000e+00, // 251
 0.000000000000000e+00, // 252
 0.000000000000000e+00, // 253
 0.000000000000000e+00, // 254
 0.000000000000000e+00, // 255
 0.000000000000000e+00, // 256
 0.000000000000000e+00, // 257
 0.000000000000000e+00, // 258
 0.000000000000000e+00, // 259
 0.000000000000000e+00, // 260
 0.000000000000000e+00, // 261
 0.000000000000000e+00, // 262
 0.000000000000000e+00, // 263
 0.000000000000000e+00, // 264
 0.000000000000000e+00, // 265
 0.000000000000000e+00, // 266
 0.000000000000000e+00, // 267
 0.000000000000000e+00, // 268
 0.000000000000000e+00, // 269
 0.000000000000000e+00, // 270
 0.000000000000000e+00, // 271
 0.000000000000000e+00, // 272
 0.000000000000000e+00, // 273
 0.000000000000000e+00, // 274
 0.000000000000000e+00, // 275
 0.000000000000000e+00, // 276
 0.000000000000000e+00, // 277
 0.000000000000000e+00, // 278
 0.000000000000000e+00, // 279
 0.000000000000000e+00, // 280
 0.000000000000000e+00, // 281
 0.000000000000000e+00, // 282
 0.000000000000000e+00, // 283
 0.000000000000000e+00, // 284
 0.000000000000000e+00, // 285
 0.000000000000000e+00, // 286
 0.000000000000000e+00, // 287
 0.000000000000000e+00, // 288
 0.000000000000000e+00, // 289
 0.000000000000000e+00, // 290
 0.000000000000000e+00, // 291
 0.000000000000000e+00, // 292
 0.000000000000000e+00, // 293
 0.000000000000000e+00, // 294
 0.000000000000000e+00, // 295
 0.000000000000000e+00, // 296
 0.000000000000000e+00, // 297
 0.000000000000000e+00, // 298
 0.000000000000000e+00, // 299
 0.000000000000000e+00, // 300
 0.000000000000000e+00, // 301
 0.000000000000000e+00, // 302
 0.000000000000000e+00, // 303
 0.000000000000000e+00, // 304
 0.000000000000000e+00, // 305
 0.000000000000000e+00, // 306
 0.000000000000000e+00, // 307
 0.000000000000000e+00, // 308
 0.000000000000000e+00, // 309
 0.000000000000000e+00, // 310
 0.000000000000000e+00, // 311
 0.000000000000000e+00, // 312
 0.000000000000000e+00, // 313
 0.000000000000000e+00, // 314
 0.000000000000000e+00, // 315
 0.000000000000000e+00, // 316
 0.000000000000000e+00, // 317
 0.000000000000000e+00, // 318
 0.000000000000000e+00, // 319
 0.000000000000000e+00, // 320
 0.000000000000000e+00, // 321
 0.000000000000000e+00, // 322
 0.000000000000000e+00, // 323
 0.000000000000000e+00, // 324
 0.000000000000000e+00, // 325
 0.000000000000000e+00, // 326
 0.000000000000000e+00, // 327
 0.000000000000000e+00, // 328
 0.000000000000000e+00, // 329
 0.000000000000000e+00, // 330
 0.000000000000000e+00, // 331
 0.000000000000000e+00, // 332
 0.000000000000000e+00, // 333
 0.000000000000000e+00, // 334
 0.000000000000000e+00, // 335
 0.000000000000000e+00, // 336
 0.000000000000000e+00, // 337
 0.000000000000000e+00, // 338
 0.000000000000000e+00, // 339
 0.000000000000000e+00, // 340
 0.000000000000000e+00, // 341
 0.000000000000000e+00, // 342
 0.000000000000000e+00, // 343
 0.000000000000000e+00, // 344
 0.000000000000000e+00, // 345
 0.000000000000000e+00, // 346
 0.000000000000000e+00, // 347
 0.000000000000000e+00, // 348
 0.000000000000000e+00, // 349
 0.000000000000000e+00, // 350
 0.000000000000000e+00, // 351
 0.000000000000000e+00, // 352
 0.000000000000000e+00, // 353
 0.000000000000000e+00, // 354
 0.000000000000000e+00, // 355
 0.000000000000000e+00, // 356
 0.000000000000000e+00, // 357
 0.000000000000000e+00, // 358
 0.000000000000000e+00, // 359
 0.000000000000000e+00, // 360
 0.000000000000000e+00, // 361
 0.000000000000000e+00, // 362
 0.000000000000000e+00, // 363
 0.000000000000000e+00, // 364
 0.000000000000000e+00, // 365
 0.000000000000000e+00, // 366
 0.000000000000000e+00, // 367
 0.000000000000000e+00, // 368
 0.000000000000000e+00, // 369
 0.000000000000000e+00, // 370
 0.000000000000000e+00, // 371
 0.000000000000000e+00, // 372
 0.000000000000000e+00, // 373
 0.000000000000000e+00, // 374
 0.000000000000000e+00, // 375
 0.000000000000000e+00, // 376
 0.000000000000000e+00, // 377
 0.000000000000000e+00, // 378
 0.000000000000000e+00, // 379
 0.000000000000000e+00, // 380
 0.000000000000000e+00, // 381
 0.000000000000000e+00, // 382
 0.000000000000000e+00, // 383
 0.000000000000000e+00, // 384
 0.000000000000000e+00, // 385
 0.000000000000000e+00, // 386
 0.000000000000000e+00, // 387
 0.000000000000000e+00, // 388
 0.000000000000000e+00, // 389
 0.000000000000000e+00, // 390
 0.000000000000000e+00, // 391
 0.000000000000000e+00, // 392
 0.000000000000000e+00, // 393
 0.000000000000000e+00, // 394
 0.000000000000000e+00, // 395
 0.000000000000000e+00, // 396
 0.000000000000000e+00, // 397
 0.000000000000000e+00, // 398
 0.000000000000000e+00, // 399
 0.000000000000000e+00, // 400
 0.000000000000000e+00, // 401
 0.000000000000000e+00, // 402
 0.000000000000000e+00, // 403
 0.000000000000000e+00, // 404
 0.000000000000000e+00, // 405
 0.000000000000000e+00, // 406
 0.000000000000000e+00, // 407
 0.000000000000000e+00, // 408
 0.000000000000000e+00, // 409
 0.000000000000000e+00, // 410
 0.000000000000000e+00, // 411
 0.000000000000000e+00, // 412
 0.000000000000000e+00, // 413
 0.000000000000000e+00, // 414
 0.000000000000000e+00, // 415
 0.000000000000000e+00, // 416
 0.000000000000000e+00, // 417
 0.000000000000000e+00, // 418
 0.000000000000000e+00, // 419
 0.000000000000000e+00, // 420
 0.000000000000000e+00, // 421
 0.000000000000000e+00, // 422
 0.000000000000000e+00, // 423
 0.000000000000000e+00, // 424
 0.000000000000000e+00, // 425
 0.000000000000000e+00, // 426
 0.000000000000000e+00, // 427
 0.000000000000000e+00, // 428
 0.000000000000000e+00, // 429
 0.000000000000000e+00, // 430
 0.000000000000000e+00, // 431
 0.000000000000000e+00, // 432
 0.000000000000000e+00, // 433
 0.000000000000000e+00, // 434
 0.000000000000000e+00, // 435
 0.000000000000000e+00, // 436
 0.000000000000000e+00, // 437
 0.000000000000000e+00, // 438
 0.000000000000000e+00, // 439
 0.000000000000000e+00, // 440
 0.000000000000000e+00, // 441
 0.000000000000000e+00, // 442
 0.000000000000000e+00, // 443
 0.000000000000000e+00, // 444
 0.000000000000000e+00, // 445
 0.000000000000000e+00, // 446
 0.000000000000000e+00, // 447
 0.000000000000000e+00, // 448
 0.000000000000000e+00, // 449
 0.000000000000000e+00, // 450
 0.000000000000000e+00, // 451
 0.000000000000000e+00, // 452
 0.000000000000000e+00, // 453
 0.000000000000000e+00, // 454
 0.000000000000000e+00, // 455
 0.000000000000000e+00, // 456
 0.000000000000000e+00, // 457
 0.000000000000000e+00, // 458
 0.000000000000000e+00, // 459
 0.000000000000000e+00, // 460
 0.000000000000000e+00, // 461
 0.000000000000000e+00, // 462
 0.000000000000000e+00, // 463
 0.000000000000000e+00, // 464
 0.000000000000000e+00, // 465
 0.000000000000000e+00, // 466
 0.000000000000000e+00, // 467
 0.000000000000000e+00, // 468
 0.000000000000000e+00, // 469
 0.000000000000000e+00, // 470
 0.000000000000000e+00, // 471
 0.000000000000000e+00, // 472
 0.000000000000000e+00, // 473
 0.000000000000000e+00, // 474
 0.000000000000000e+00, // 475
 0.000000000000000e+00, // 476
 0.000000000000000e+00, // 477
 0.000000000000000e+00, // 478
 0.000000000000000e+00, // 479
 0.000000000000000e+00, // 480
 0.000000000000000e+00, // 481
 0.000000000000000e+00, // 482
 0.000000000000000e+00, // 483
 0.000000000000000e+00, // 484
 0.000000000000000e+00, // 485
 0.000000000000000e+00, // 486
 0.000000000000000e+00, // 487
 0.000000000000000e+00, // 488
 0.000000000000000e+00, // 489
 0.000000000000000e+00, // 490
 0.000000000000000e+00, // 491
 0.000000000000000e+00, // 492
 0.000000000000000e+00, // 493
 0.000000000000000e+00, // 494
 0.000000000000000e+00, // 495
 0.000000000000000e+00, // 496
 0.000000000000000e+00, // 497
 0.000000000000000e+00, // 498
 0.000000000000000e+00, // 499
 0.000000000000000e+00, // 500
 0.000000000000000e+00, // 501
 0.000000000000000e+00, // 502
 0.000000000000000e+00, // 503
 0.000000000000000e+00, // 504
 0.000000000000000e+00, // 505
 0.000000000000000e+00, // 506
 0.000000000000000e+00, // 507
 0.000000000000000e+00, // 508
 0.000000000000000e+00, // 509
 0.000000000000000e+00, // 510
 0.000000000000000e+00, // 511
 0.000000000000000e+00, // 512
 0.000000000000000e+00, // 513
 0.000000000000000e+00, // 514
 0.000000000000000e+00, // 515
 0.000000000000000e+00, // 516
 0.000000000000000e+00, // 517
 0.000000000000000e+00, // 518
 0.000000000000000e+00, // 519
 0.000000000000000e+00, // 520
 0.000000000000000e+00, // 521
 0.000000000000000e+00, // 522
 0.000000000000000e+00, // 523
 0.000000000000000e+00, // 524
 0.000000000000000e+00, // 525
 0.000000000000000e+00, // 526
 0.000000000000000e+00, // 527
 0.000000000000000e+00, // 528
 0.000000000000000e+00, // 529
 0.000000000000000e+00, // 530
 0.000000000000000e+00, // 531
 0.000000000000000e+00, // 532
 0.000000000000000e+00, // 533
 0.000000000000000e+00, // 534
 0.000000000000000e+00, // 535
 0.000000000000000e+00, // 536
 0.000000000000000e+00, // 537
 0.000000000000000e+00, // 538
 0.000000000000000e+00, // 539
 0.000000000000000e+00, // 540
 0.000000000000000e+00, // 541
 0.000000000000000e+00, // 542
 0.000000000000000e+00, // 543
 0.000000000000000e+00, // 544
 0.000000000000000e+00, // 545
 0.000000000000000e+00, // 546
 0.000000000000000e+00, // 547
 0.000000000000000e+00, // 548
 0.000000000000000e+00, // 549
 0.000000000000000e+00, // 550
 0.000000000000000e+00, // 551
 0.000000000000000e+00, // 552
 0.000000000000000e+00, // 553
 0.000000000000000e+00, // 554
 0.000000000000000e+00, // 555
 0.000000000000000e+00, // 556
 0.000000000000000e+00, // 557
 0.000000000000000e+00, // 558
 0.000000000000000e+00, // 559
 0.000000000000000e+00, // 560
 0.000000000000000e+00, // 561
 0.000000000000000e+00, // 562
 0.000000000000000e+00, // 563
 0.000000000000000e+00, // 564
 0.000000000000000e+00, // 565
 0.000000000000000e+00, // 566
 0.000000000000000e+00, // 567
 0.000000000000000e+00, // 568
 0.000000000000000e+00, // 569
 0.000000000000000e+00, // 570
 0.000000000000000e+00, // 571
 0.000000000000000e+00, // 572
 0.000000000000000e+00, // 573
 0.000000000000000e+00, // 574
 0.000000000000000e+00, // 575
 0.000000000000000e+00, // 576
 0.000000000000000e+00, // 577
 0.000000000000000e+00, // 578
 0.000000000000000e+00, // 579
 0.000000000000000e+00, // 580
 0.000000000000000e+00, // 581
 0.000000000000000e+00, // 582
 0.000000000000000e+00, // 583
 0.000000000000000e+00, // 584
 0.000000000000000e+00, // 585
 0.000000000000000e+00, // 586
 0.000000000000000e+00, // 587
 0.000000000000000e+00, // 588
 0.000000000000000e+00, // 589
 0.000000000000000e+00, // 590
 0.000000000000000e+00, // 591
 0.000000000000000e+00, // 592
 0.000000000000000e+00, // 593
 0.000000000000000e+00, // 594
 0.000000000000000e+00, // 595
 0.000000000000000e+00, // 596
 0.000000000000000e+00, // 597
 0.000000000000000e+00, // 598
 0.000000000000000e+00, // 599
 0.000000000000000e+00, // 600
 0.000000000000000e+00, // 601
 0.000000000000000e+00, // 602
 0.000000000000000e+00, // 603
 0.000000000000000e+00, // 604
 0.000000000000000e+00, // 605
 0.000000000000000e+00, // 606
 0.000000000000000e+00, // 607
 0.000000000000000e+00, // 608
 0.000000000000000e+00, // 609
 0.000000000000000e+00, // 610
 0.000000000000000e+00, // 611
 0.000000000000000e+00, // 612
 0.000000000000000e+00, // 613
 0.000000000000000e+00, // 614
 0.000000000000000e+00, // 615
 0.000000000000000e+00, // 616
 0.000000000000000e+00, // 617
 0.000000000000000e+00, // 618
 0.000000000000000e+00, // 619
 0.000000000000000e+00, // 620
 0.000000000000000e+00, // 621
 0.000000000000000e+00, // 622
 0.000000000000000e+00, // 623
 0.000000000000000e+00, // 624
 0.000000000000000e+00, // 625
 0.000000000000000e+00, // 626
 0.000000000000000e+00, // 627
 0.000000000000000e+00, // 628
 0.000000000000000e+00, // 629
 0.000000000000000e+00, // 630
 0.000000000000000e+00, // 631
 0.000000000000000e+00, // 632
 0.000000000000000e+00, // 633
 0.000000000000000e+00, // 634
 0.000000000000000e+00, // 635
 0.000000000000000e+00, // 636
 0.000000000000000e+00, // 637
 0.000000000000000e+00, // 638
 0.000000000000000e+00, // 639
 0.000000000000000e+00, // 640
 0.000000000000000e+00, // 641
 0.000000000000000e+00, // 642
 0.000000000000000e+00, // 643
 0.000000000000000e+00, // 644
 0.000000000000000e+00, // 645
 0.000000000000000e+00, // 646
 0.000000000000000e+00, // 647
 0.000000000000000e+00, // 648
 0.000000000000000e+00, // 649
 0.000000000000000e+00, // 650
 0.000000000000000e+00, // 651
 0.000000000000000e+00, // 652
 0.000000000000000e+00, // 653
 0.000000000000000e+00, // 654
 0.000000000000000e+00, // 655
 0.000000000000000e+00, // 656
 0.000000000000000e+00, // 657
 0.000000000000000e+00, // 658
 0.000000000000000e+00, // 659
 0.000000000000000e+00, // 660
 0.000000000000000e+00, // 661
 0.000000000000000e+00, // 662
 0.000000000000000e+00, // 663
 0.000000000000000e+00, // 664
 0.000000000000000e+00, // 665
 0.000000000000000e+00, // 666
 0.000000000000000e+00, // 667
 0.000000000000000e+00, // 668
 0.000000000000000e+00, // 669
 0.000000000000000e+00, // 670
 0.000000000000000e+00, // 671
 0.000000000000000e+00, // 672
 0.000000000000000e+00, // 673
 0.000000000000000e+00, // 674
 0.000000000000000e+00, // 675
 0.000000000000000e+00, // 676
 0.000000000000000e+00, // 677
 0.000000000000000e+00, // 678
 0.000000000000000e+00, // 679
 0.000000000000000e+00, // 680
 0.000000000000000e+00, // 681
 0.000000000000000e+00, // 682
 0.000000000000000e+00, // 683
 0.000000000000000e+00, // 684
 0.000000000000000e+00, // 685
 0.000000000000000e+00, // 686
 0.000000000000000e+00, // 687
 0.000000000000000e+00, // 688
 0.000000000000000e+00, // 689
 0.000000000000000e+00, // 690
 0.000000000000000e+00, // 691
 0.000000000000000e+00, // 692
 0.000000000000000e+00, // 693
 0.000000000000000e+00, // 694
 0.000000000000000e+00, // 695
 0.000000000000000e+00, // 696
 0.000000000000000e+00, // 697
 0.000000000000000e+00, // 698
 0.000000000000000e+00, // 699
 0.000000000000000e+00, // 700
 0.000000000000000e+00, // 701
 0.000000000000000e+00, // 702
 0.000000000000000e+00, // 703
 0.000000000000000e+00, // 704
 0.000000000000000e+00, // 705
 0.000000000000000e+00, // 706
 0.000000000000000e+00, // 707
 0.000000000000000e+00, // 708
 0.000000000000000e+00, // 709
 0.000000000000000e+00, // 710
 0.000000000000000e+00, // 711
 0.000000000000000e+00, // 712
 0.000000000000000e+00, // 713
 0.000000000000000e+00, // 714
 0.000000000000000e+00, // 715
 0.000000000000000e+00, // 716
 0.000000000000000e+00, // 717
 0.000000000000000e+00, // 718
 0.000000000000000e+00, // 719
 0.000000000000000e+00, // 720
 0.000000000000000e+00, // 721
 0.000000000000000e+00, // 722
 0.000000000000000e+00, // 723
 0.000000000000000e+00, // 724
 0.000000000000000e+00, // 725
 0.000000000000000e+00, // 726
 0.000000000000000e+00, // 727
 0.000000000000000e+00, // 728
 0.000000000000000e+00, // 729
 0.000000000000000e+00, // 730
 0.000000000000000e+00, // 731
 0.000000000000000e+00, // 732
 0.000000000000000e+00, // 733
 0.000000000000000e+00, // 734
 0.000000000000000e+00, // 735
 0.000000000000000e+00, // 736
 0.000000000000000e+00, // 737
 0.000000000000000e+00, // 738
 0.000000000000000e+00, // 739
 0.000000000000000e+00, // 740
 0.000000000000000e+00, // 741
 0.000000000000000e+00, // 742
 0.000000000000000e+00, // 743
 0.000000000000000e+00, // 744
 0.000000000000000e+00, // 745
 0.000000000000000e+00, // 746
 0.000000000000000e+00, // 747
 0.000000000000000e+00, // 748
 0.000000000000000e+00, // 749
 0.000000000000000e+00, // 750
 0.000000000000000e+00, // 751
 0.000000000000000e+00, // 752
 0.000000000000000e+00, // 753
 0.000000000000000e+00, // 754
 0.000000000000000e+00, // 755
 0.000000000000000e+00, // 756
 0.000000000000000e+00, // 757
 0.000000000000000e+00, // 758
 0.000000000000000e+00, // 759
 0.000000000000000e+00, // 760
 0.000000000000000e+00, // 761
 0.000000000000000e+00, // 762
 0.000000000000000e+00, // 763
 0.000000000000000e+00, // 764
 0.000000000000000e+00, // 765
 0.000000000000000e+00, // 766
 0.000000000000000e+00, // 767
 0.000000000000000e+00, // 768
 0.000000000000000e+00, // 769
 0.000000000000000e+00, // 770
 0.000000000000000e+00, // 771
 0.000000000000000e+00, // 772
 0.000000000000000e+00, // 773
 0.000000000000000e+00, // 774
 0.000000000000000e+00, // 775
 0.000000000000000e+00, // 776
 0.000000000000000e+00, // 777
 0.000000000000000e+00, // 778
 0.000000000000000e+00, // 779
 0.000000000000000e+00, // 780
 0.000000000000000e+00, // 781
 0.000000000000000e+00, // 782
 0.000000000000000e+00, // 783
 0.000000000000000e+00, // 784
 0.000000000000000e+00, // 785
 0.000000000000000e+00, // 786
 0.000000000000000e+00, // 787
 0.000000000000000e+00, // 788
 0.000000000000000e+00, // 789
 0.000000000000000e+00, // 790
 0.000000000000000e+00, // 791
 0.000000000000000e+00, // 792
 0.000000000000000e+00, // 793
 0.000000000000000e+00, // 794
 0.000000000000000e+00, // 795
 0.000000000000000e+00, // 796
 0.000000000000000e+00, // 797
 0.000000000000000e+00, // 798
 0.000000000000000e+00, // 799
 0.000000000000000e+00, // 800
 0.000000000000000e+00, // 801
 0.000000000000000e+00, // 802
 0.000000000000000e+00, // 803
 0.000000000000000e+00, // 804
 0.000000000000000e+00, // 805
 0.000000000000000e+00, // 806
 0.000000000000000e+00, // 807
 0.000000000000000e+00, // 808
 0.000000000000000e+00, // 809
 0.000000000000000e+00, // 810
 0.000000000000000e+00, // 811
 0.000000000000000e+00, // 812
 0.000000000000000e+00, // 813
 0.000000000000000e+00, // 814
 0.000000000000000e+00, // 815
 0.000000000000000e+00, // 816
 0.000000000000000e+00, // 817
 0.000000000000000e+00, // 818
 0.000000000000000e+00, // 819
 0.000000000000000e+00, // 820
 0.000000000000000e+00, // 821
 0.000000000000000e+00, // 822
 0.000000000000000e+00, // 823
 0.000000000000000e+00, // 824
 0.000000000000000e+00, // 825
 0.000000000000000e+00, // 826
 0.000000000000000e+00, // 827
 0.000000000000000e+00, // 828
 0.000000000000000e+00, // 829
 0.000000000000000e+00, // 830
 0.000000000000000e+00, // 831
 0.000000000000000e+00, // 832
 0.000000000000000e+00, // 833
 0.000000000000000e+00, // 834
 0.000000000000000e+00, // 835
 0.000000000000000e+00, // 836
 0.000000000000000e+00, // 837
 0.000000000000000e+00, // 838
 0.000000000000000e+00, // 839
 0.000000000000000e+00, // 840
 0.000000000000000e+00, // 841
 0.000000000000000e+00, // 842
 0.000000000000000e+00, // 843
 0.000000000000000e+00, // 844
 0.000000000000000e+00, // 845
 0.000000000000000e+00, // 846
 0.000000000000000e+00, // 847
 0.000000000000000e+00, // 848
 0.000000000000000e+00, // 849
 0.000000000000000e+00, // 850
 0.000000000000000e+00, // 851
 0.000000000000000e+00, // 852
 0.000000000000000e+00, // 853
 0.000000000000000e+00, // 854
 0.000000000000000e+00, // 855
 0.000000000000000e+00, // 856
 0.000000000000000e+00, // 857
 0.000000000000000e+00, // 858
 0.000000000000000e+00, // 859
 0.000000000000000e+00, // 860
 0.000000000000000e+00, // 861
 0.000000000000000e+00, // 862
 0.000000000000000e+00, // 863
 0.000000000000000e+00, // 864
 0.000000000000000e+00, // 865
 0.000000000000000e+00, // 866
 0.000000000000000e+00, // 867
 0.000000000000000e+00, // 868
 0.000000000000000e+00, // 869
 0.000000000000000e+00, // 870
 0.000000000000000e+00, // 871
 0.000000000000000e+00, // 872
 0.000000000000000e+00, // 873
 0.000000000000000e+00, // 874
 0.000000000000000e+00, // 875
 0.000000000000000e+00, // 876
 0.000000000000000e+00, // 877
 0.000000000000000e+00, // 878
 0.000000000000000e+00, // 879
 0.000000000000000e+00, // 880
 0.000000000000000e+00, // 881
 0.000000000000000e+00, // 882
 0.000000000000000e+00, // 883
 0.000000000000000e+00, // 884
 0.000000000000000e+00, // 885
 0.000000000000000e+00, // 886
 0.000000000000000e+00, // 887
 0.000000000000000e+00, // 888
 0.000000000000000e+00, // 889
 0.000000000000000e+00, // 890
 0.000000000000000e+00, // 891
 0.000000000000000e+00, // 892
 0.000000000000000e+00, // 893
 0.000000000000000e+00, // 894
 0.000000000000000e+00, // 895
 0.000000000000000e+00, // 896
 0.000000000000000e+00, // 897
 0.000000000000000e+00, // 898
 0.000000000000000e+00, // 899
 0.000000000000000e+00, // 900
 0.000000000000000e+00, // 901
 0.000000000000000e+00, // 902
 0.000000000000000e+00, // 903
 0.000000000000000e+00, // 904
 0.000000000000000e+00, // 905
 0.000000000000000e+00, // 906
 0.000000000000000e+00, // 907
 0.000000000000000e+00, // 908
 0.000000000000000e+00, // 909
 0.000000000000000e+00, // 910
 0.000000000000000e+00, // 911
 0.000000000000000e+00, // 912
 0.000000000000000e+00, // 913
 0.000000000000000e+00, // 914
 0.000000000000000e+00, // 915
 0.000000000000000e+00, // 916
 0.000000000000000e+00, // 917
 0.000000000000000e+00, // 918
 0.000000000000000e+00, // 919
 0.000000000000000e+00, // 920
 0.000000000000000e+00, // 921
 0.000000000000000e+00, // 922
 0.000000000000000e+00, // 923
 0.000000000000000e+00, // 924
 0.000000000000000e+00, // 925
 0.000000000000000e+00, // 926
 0.000000000000000e+00, // 927
 0.000000000000000e+00, // 928
 0.000000000000000e+00, // 929
 0.000000000000000e+00, // 930
 0.000000000000000e+00, // 931
 0.000000000000000e+00, // 932
 0.000000000000000e+00, // 933
 0.000000000000000e+00, // 934
 0.000000000000000e+00, // 935
 0.000000000000000e+00, // 936
 0.000000000000000e+00, // 937
 0.000000000000000e+00, // 938
 0.000000000000000e+00, // 939
 0.000000000000000e+00, // 940
 0.000000000000000e+00, // 941
 0.000000000000000e+00, // 942
 0.000000000000000e+00, // 943
 0.000000000000000e+00, // 944
 0.000000000000000e+00, // 945
 0.000000000000000e+00, // 946
 0.000000000000000e+00, // 947
 0.000000000000000e+00, // 948
 0.000000000000000e+00, // 949
 0.000000000000000e+00, // 950
 0.000000000000000e+00, // 951
 0.000000000000000e+00, // 952
 0.000000000000000e+00, // 953
 0.000000000000000e+00, // 954
 0.000000000000000e+00, // 955
 0.000000000000000e+00, // 956
 0.000000000000000e+00, // 957
 0.000000000000000e+00, // 958
 0.000000000000000e+00, // 959
 0.000000000000000e+00, // 960
 0.000000000000000e+00, // 961
 0.000000000000000e+00, // 962
 0.000000000000000e+00, // 963
 0.000000000000000e+00, // 964
 0.000000000000000e+00, // 965
 0.000000000000000e+00, // 966
 0.000000000000000e+00, // 967
 0.000000000000000e+00, // 968
 0.000000000000000e+00, // 969
 0.000000000000000e+00, // 970
 0.000000000000000e+00, // 971
 0.000000000000000e+00, // 972
 0.000000000000000e+00, // 973
 0.000000000000000e+00, // 974
 0.000000000000000e+00, // 975
 0.000000000000000e+00, // 976
 0.000000000000000e+00, // 977
 0.000000000000000e+00, // 978
 0.000000000000000e+00, // 979
 0.000000000000000e+00, // 980
 0.000000000000000e+00, // 981
 0.000000000000000e+00, // 982
 0.000000000000000e+00, // 983
 0.000000000000000e+00, // 984
 0.000000000000000e+00, // 985
 0.000000000000000e+00, // 986
 0.000000000000000e+00, // 987
 0.000000000000000e+00, // 988
 0.000000000000000e+00, // 989
 0.000000000000000e+00, // 990
 0.000000000000000e+00, // 991
 0.000000000000000e+00, // 992
 0.000000000000000e+00, // 993
 0.000000000000000e+00, // 994
 0.000000000000000e+00, // 995
 0.000000000000000e+00, // 996
 0.000000000000000e+00, // 997
 0.000000000000000e+00, // 998
 0.000000000000000e+00, // 999
 0.000000000000000e+00, // 1000
 0.000000000000000e+00, // 1001
 0.000000000000000e+00, // 1002
 0.000000000000000e+00, // 1003
 0.000000000000000e+00, // 1004
 0.000000000000000e+00, // 1005
 0.000000000000000e+00, // 1006
 0.000000000000000e+00, // 1007
 0.000000000000000e+00, // 1008
 0.000000000000000e+00, // 1009
 0.000000000000000e+00, // 1010
 0.000000000000000e+00, // 1011
 0.000000000000000e+00, // 1012
 0.000000000000000e+00, // 1013
 0.000000000000000e+00, // 1014
 0.000000000000000e+00, // 1015
 0.000000000000000e+00, // 1016
 0.000000000000000e+00, // 1017
 0.000000000000000e+00, // 1018
 0.000000000000000e+00, // 1019
 0.000000000000000e+00, // 1020
 0.000000000000000e+00, // 1021
 0.000000000000000e+00, // 1022
 0.000000000000000e+00, // 1023
 0.000000000000000e+00, // 1024
 0.000000000000000e+00, // 1025
 0.000000000000000e+00, // 1026
 0.000000000000000e+00, // 1027
 0.000000000000000e+00, // 1028
 0.000000000000000e+00, // 1029
 0.000000000000000e+00, // 1030
 0.000000000000000e+00, // 1031
 0.000000000000000e+00, // 1032
 0.000000000000000e+00, // 1033
 0.000000000000000e+00, // 1034
 0.000000000000000e+00, // 1035
 0.000000000000000e+00, // 1036
 0.000000000000000e+00, // 1037
 0.000000000000000e+00, // 1038
 0.000000000000000e+00, // 1039
 0.000000000000000e+00, // 1040
 0.000000000000000e+00, // 1041
 0.000000000000000e+00, // 1042
 0.000000000000000e+00, // 1043
 0.000000000000000e+00, // 1044
 0.000000000000000e+00, // 1045
 0.000000000000000e+00, // 1046
 0.000000000000000e+00, // 1047
 0.000000000000000e+00, // 1048
 0.000000000000000e+00, // 1049
 0.000000000000000e+00, // 1050
 0.000000000000000e+00, // 1051
 0.000000000000000e+00, // 1052
 0.000000000000000e+00, // 1053
 0.000000000000000e+00, // 1054
 0.000000000000000e+00, // 1055
 0.000000000000000e+00, // 1056
 0.000000000000000e+00, // 1057
 0.000000000000000e+00, // 1058
 0.000000000000000e+00, // 1059
 0.000000000000000e+00, // 1060
 0.000000000000000e+00, // 1061
 0.000000000000000e+00, // 1062
 0.000000000000000e+00, // 1063
 0.000000000000000e+00, // 1064
 0.000000000000000e+00, // 1065
 0.000000000000000e+00, // 1066
 0.000000000000000e+00, // 1067
 0.000000000000000e+00, // 1068
 0.000000000000000e+00, // 1069
 0.000000000000000e+00, // 1070
 0.000000000000000e+00, // 1071
 0.000000000000000e+00, // 1072
 0.000000000000000e+00, // 1073
 0.000000000000000e+00, // 1074
 0.000000000000000e+00, // 1075
 0.000000000000000e+00, // 1076
 0.000000000000000e+00, // 1077
 0.000000000000000e+00, // 1078
 0.000000000000000e+00, // 1079
 0.000000000000000e+00, // 1080
 0.000000000000000e+00, // 1081
 0.000000000000000e+00, // 1082
 0.000000000000000e+00, // 1083
 0.000000000000000e+00, // 1084
 0.000000000000000e+00, // 1085
 0.000000000000000e+00, // 1086
 0.000000000000000e+00, // 1087
 0.000000000000000e+00, // 1088
 0.000000000000000e+00, // 1089
 0.000000000000000e+00, // 1090
 0.000000000000000e+00, // 1091
 0.000000000000000e+00, // 1092
 0.000000000000000e+00, // 1093
 0.000000000000000e+00, // 1094
 0.000000000000000e+00, // 1095
 0.000000000000000e+00, // 1096
 0.000000000000000e+00, // 1097
 0.000000000000000e+00, // 1098
 0.000000000000000e+00, // 1099
 0.000000000000000e+00, // 1100
 0.000000000000000e+00, // 1101
 0.000000000000000e+00, // 1102
 0.000000000000000e+00, // 1103
 0.000000000000000e+00, // 1104
 0.000000000000000e+00, // 1105
 0.000000000000000e+00, // 1106
 0.000000000000000e+00, // 1107
 0.000000000000000e+00, // 1108
 0.000000000000000e+00, // 1109
 0.000000000000000e+00, // 1110
 0.000000000000000e+00, // 1111
 0.000000000000000e+00, // 1112
 0.000000000000000e+00, // 1113
 0.000000000000000e+00, // 1114
 0.000000000000000e+00, // 1115
 0.000000000000000e+00, // 1116
 0.000000000000000e+00, // 1117
 0.000000000000000e+00, // 1118
 0.000000000000000e+00, // 1119
 0.000000000000000e+00, // 1120
 0.000000000000000e+00, // 1121
 0.000000000000000e+00, // 1122
 0.000000000000000e+00, // 1123
 0.000000000000000e+00, // 1124
 0.000000000000000e+00, // 1125
 0.000000000000000e+00, // 1126
 0.000000000000000e+00, // 1127
 0.000000000000000e+00, // 1128
 0.000000000000000e+00, // 1129
 0.000000000000000e+00, // 1130
 0.000000000000000e+00, // 1131
 0.000000000000000e+00, // 1132
 0.000000000000000e+00, // 1133
 0.000000000000000e+00, // 1134
 0.000000000000000e+00, // 1135
 0.000000000000000e+00, // 1136
 0.000000000000000e+00, // 1137
 0.000000000000000e+00, // 1138
 0.000000000000000e+00, // 1139
 0.000000000000000e+00, // 1140
 0.000000000000000e+00, // 1141
 0.000000000000000e+00, // 1142
 0.000000000000000e+00, // 1143
 0.000000000000000e+00, // 1144
 0.000000000000000e+00, // 1145
 0.000000000000000e+00, // 1146
 0.000000000000000e+00, // 1147
 0.000000000000000e+00, // 1148
 0.000000000000000e+00, // 1149
 0.000000000000000e+00, // 1150
 0.000000000000000e+00, // 1151
 0.000000000000000e+00, // 1152
 0.000000000000000e+00, // 1153
 0.000000000000000e+00, // 1154
 0.000000000000000e+00, // 1155
 0.000000000000000e+00, // 1156
 0.000000000000000e+00, // 1157
 0.000000000000000e+00, // 1158
 0.000000000000000e+00, // 1159
 0.000000000000000e+00, // 1160
 0.000000000000000e+00, // 1161
 0.000000000000000e+00, // 1162
 0.000000000000000e+00, // 1163
 0.000000000000000e+00, // 1164
 0.000000000000000e+00, // 1165
 0.000000000000000e+00, // 1166
 0.000000000000000e+00, // 1167
 0.000000000000000e+00, // 1168
 0.000000000000000e+00, // 1169
 0.000000000000000e+00, // 1170
 0.000000000000000e+00, // 1171
 0.000000000000000e+00, // 1172
 0.000000000000000e+00, // 1173
 0.000000000000000e+00, // 1174
 0.000000000000000e+00, // 1175
 0.000000000000000e+00, // 1176
 0.000000000000000e+00, // 1177
 0.000000000000000e+00, // 1178
 0.000000000000000e+00, // 1179
 0.000000000000000e+00, // 1180
 0.000000000000000e+00, // 1181
 0.000000000000000e+00; // 1182

}
